////Main Module For Processing
module LeNet1 (clk, rst, data, answer, result);
  input clk, rst;
  input [784*16 - 1:0] data;
  input [9:0] answer;
  output reg result;
  
  wire [576*16 - 1:0] data_11, data_12, data_13, data_14;
  
  //Parameters
  parameter CONV1_WEIGHTS_ROW = 4,
    CONV1_WEIGHTS_COLUMN = 25,
    CONV1_BIAS_ROW = 4,
    CONV2_WEIGHTS_ROW = 12,
    CONV2_WEIGHTS_COLUMN = 100,
    CONV2_BIAS_ROW = 12,
    FC1_WEIGHTS_ROW = 10,
    FC1_WEIGHTS_COLUMN = 192,
    FC1_BIAS_ROW = 10,
    FP_LENGTH = 16;
    
    
  //Memory arrays in which all the parameters will be imported
  reg [FP_LENGTH - 1:0] CONV1_WEIGHTS_M [CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1:0];
  reg [FP_LENGTH - 1:0] CONV1_BIAS_M [CONV1_BIAS_ROW - 1:0];
  reg [FP_LENGTH - 1:0] CONV2_WEIGHTS_M [CONV2_WEIGHTS_ROW*CONV2_WEIGHTS_COLUMN - 1:0];
  reg [FP_LENGTH - 1:0] CONV2_BIAS_M [CONV2_BIAS_ROW - 1:0];
  reg [FP_LENGTH - 1:0] FC1_WEIGHTS_M [FC1_WEIGHTS_ROW*FC1_WEIGHTS_COLUMN - 1:0];
  reg [FP_LENGTH - 1:0] FC1_BIAS_M [FC1_BIAS_ROW - 1:0];
  
  initial begin
   //Importing all required files in memory arrays
   $readmemb("C:/Users/king/Documents/Jupyter/HA/Files/conv1_weight.txt", CONV1_WEIGHTS_M);
   $readmemb("C:/Users/king/Documents/Jupyter/HA/Files/conv1_bias.txt", CONV1_BIAS_M);
   $readmemb("C:/Users/king/Documents/Jupyter/HA/Files/conv2_weight.txt", CONV2_WEIGHTS_M);
   $readmemb("C:/Users/king/Documents/Jupyter/HA/Files/conv2_bias.txt", CONV2_BIAS_M);
   $readmemb("C:/Users/king/Documents/Jupyter/HA/Files/fc1_weight.txt", FC1_WEIGHTS_M);
   $readmemb("C:/Users/king/Documents/Jupyter/HA/Files/fc1_bias.txt", FC1_BIAS_M);
   //$readmemb("C:/Users/king/Documents/Jupyter/HA/Files/test_data.txt", TEST_DATA_M);
   
   
  end
  
  ////CONVOLUTION 1
  
  //FEATURE MAP 1
  Conv1_feature1 conv1_f1 (.data(data),
    .feature1Weight_0(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*0]),
    .feature1Weight_1(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*1]),
    .feature1Weight_2(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*2]),
    .feature1Weight_3(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*3]),
    .feature1Weight_4(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*4]),
    .feature1Weight_5(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*5]),
    .feature1Weight_6(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*6]),
    .feature1Weight_7(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*7]),
    .feature1Weight_8(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*8]),
    .feature1Weight_9(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*9]),
    .feature1Weight_10(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*10]),
    .feature1Weight_11(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*11]),
    .feature1Weight_12(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*12]),
    .feature1Weight_13(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*13]),
    .feature1Weight_14(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*14]),
    .feature1Weight_15(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*15]),
    .feature1Weight_16(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*16]),
    .feature1Weight_17(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*17]),
    .feature1Weight_18(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*18]),
    .feature1Weight_19(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*19]),
    .feature1Weight_20(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*20]),
    .feature1Weight_21(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*21]),
    .feature1Weight_22(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*22]),
    .feature1Weight_23(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*23]),
    .feature1Weight_24(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*24]),
    .feature1Bias(CONV1_BIAS_M [CONV1_BIAS_ROW - 1 - 1*0]),
    .data_11(data11));
    
  //FEATURE MAP 2
  Conv1_feature2 conv1_f2 (.data(data),
    .feature1Weight_0(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*25]),
    .feature1Weight_1(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*26]),
    .feature1Weight_2(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*27]),
    .feature1Weight_3(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*28]),
    .feature1Weight_4(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*29]),
    .feature1Weight_5(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*30]),
    .feature1Weight_6(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*31]),
    .feature1Weight_7(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*32]),
    .feature1Weight_8(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*33]),
    .feature1Weight_9(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*34]),
    .feature1Weight_10(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*35]),
    .feature1Weight_11(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*36]),
    .feature1Weight_12(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*37]),
    .feature1Weight_13(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*38]),
    .feature1Weight_14(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*39]),
    .feature1Weight_15(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*40]),
    .feature1Weight_16(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*41]),
    .feature1Weight_17(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*42]),
    .feature1Weight_18(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*43]),
    .feature1Weight_19(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*44]),
    .feature1Weight_20(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*45]),
    .feature1Weight_21(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*46]),
    .feature1Weight_22(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*47]),
    .feature1Weight_23(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*48]),
    .feature1Weight_24(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*49]),
    .feature1Bias(CONV1_BIAS_M [CONV1_BIAS_ROW - 1 - 1*1]),
    .data_11(data12));
    
  //FEATURE MAP 3
  Conv1_feature3 conv1_f3 (.data(data),
    .feature1Weight_0(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*50]),
    .feature1Weight_1(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*51]),
    .feature1Weight_2(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*52]),
    .feature1Weight_3(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*53]),
    .feature1Weight_4(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*54]),
    .feature1Weight_5(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*55]),
    .feature1Weight_6(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*56]),
    .feature1Weight_7(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*57]),
    .feature1Weight_8(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*58]),
    .feature1Weight_9(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*59]),
    .feature1Weight_10(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*60]),
    .feature1Weight_11(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*61]),
    .feature1Weight_12(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*62]),
    .feature1Weight_13(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*63]),
    .feature1Weight_14(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*64]),
    .feature1Weight_15(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*65]),
    .feature1Weight_16(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*66]),
    .feature1Weight_17(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*67]),
    .feature1Weight_18(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*68]),
    .feature1Weight_19(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*69]),
    .feature1Weight_20(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*70]),
    .feature1Weight_21(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*71]),
    .feature1Weight_22(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*72]),
    .feature1Weight_23(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*73]),
    .feature1Weight_24(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*74]),
    .feature1Bias(CONV1_BIAS_M [CONV1_BIAS_ROW - 1 - 1*2]),
    .data_11(data13));
    
  //FEATURE MAP 4
  Conv1_feature4 conv1_f4 (.data(data),
    .feature1Weight_0(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*75]),
    .feature1Weight_1(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*76]),
    .feature1Weight_2(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*77]),
    .feature1Weight_3(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*78]),
    .feature1Weight_4(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*79]),
    .feature1Weight_5(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*80]),
    .feature1Weight_6(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*81]),
    .feature1Weight_7(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*82]),
    .feature1Weight_8(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*83]),
    .feature1Weight_9(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*84]),
    .feature1Weight_10(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*85]),
    .feature1Weight_11(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*86]),
    .feature1Weight_12(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*87]),
    .feature1Weight_13(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*88]),
    .feature1Weight_14(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*89]),
    .feature1Weight_15(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*90]),
    .feature1Weight_16(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*91]),
    .feature1Weight_17(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*92]),
    .feature1Weight_18(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*93]),
    .feature1Weight_19(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*94]),
    .feature1Weight_20(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*95]),
    .feature1Weight_21(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*96]),
    .feature1Weight_22(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*97]),
    .feature1Weight_23(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*98]),
    .feature1Weight_24(CONV1_WEIGHTS_M[CONV1_WEIGHTS_ROW*CONV1_WEIGHTS_COLUMN - 1 - 1*99]),
    .feature1Bias(CONV1_BIAS_M [CONV1_BIAS_ROW - 1 - 1*3]),
    .data_11(data14));
    
  
  ////AVERAGE POOLING
  
  
  ////RELU
  
  
  ////COVOLUTION 2
  
  //FEATURE MAP 1
  
  //FEATURE MAP 2
  
  //FEATURE MAP 3
  
  //FEATURE MAP 4
  
  ////AVERAGE POOLING
  
  
  ////RELU
  
  
  ////FULLY CONNECTED LAYER
  
  always@ (posedge clk, negedge rst) begin
  
   if (!rst) result = 0;
   else begin
   
   end
  
  end
endmodule