//////CONVOLUTION LAYER 1

////CONVOLUTION LAYER 1 | FEATURE MAP 1
module Conv1_feature1 (
    data,
    feature1Weight_0,
    feature1Weight_1,
    feature1Weight_2,
    feature1Weight_3,
    feature1Weight_4,
    feature1Weight_5,
    feature1Weight_6,
    feature1Weight_7,
    feature1Weight_8,
    feature1Weight_9,
    feature1Weight_10,
    feature1Weight_11,
    feature1Weight_12,
    feature1Weight_13,
    feature1Weight_14,
    feature1Weight_15,
    feature1Weight_16,
    feature1Weight_17,
    feature1Weight_18,
    feature1Weight_19,
    feature1Weight_20,
    feature1Weight_21,
    feature1Weight_22,
    feature1Weight_23,
    feature1Weight_24,
    feature1Bias,
    data_11);

  parameter TEST_DATA = 784*16,
    FP_LENGTH = 16;
  input [TEST_DATA - 1:0] data;
  input [FP_LENGTH - 1:0] feature1Weight_0, feature1Weight_1, feature1Weight_2, feature1Weight_3, feature1Weight_4, feature1Weight_5, feature1Weight_6, feature1Weight_7, feature1Weight_8, feature1Weight_9, feature1Weight_10, feature1Weight_11, feature1Weight_12, feature1Weight_13, feature1Weight_14, feature1Weight_15, feature1Weight_16, feature1Weight_17, feature1Weight_18, feature1Weight_19, feature1Weight_20, feature1Weight_21, feature1Weight_22, feature1Weight_23, feature1Weight_24, feature1Bias;
  output [576*16 - 1:0] data_11;    
  
  wire [FP_LENGTH - 1:0] data_array [0:27][0:27];
  wire [FP_LENGTH - 1:0] data_11_array [0:23][0:23];
  wire [FP_LENGTH - 1:0] multi0 [0:24][0:23], multi1 [0:24][0:23], multi2 [0:24][0:23], multi3 [0:24][0:23], multi4 [0:24][0:23], multi5 [0:24][0:23], multi6 [0:24][0:23], multi7 [0:24][0:23], multi8 [0:24][0:23], multi9 [0:24][0:23], multi10 [0:24][0:23], multi11 [0:24][0:23], multi12 [0:24][0:23], multi13 [0:24][0:23], multi14 [0:24][0:23], multi15 [0:24][0:23], multi16 [0:24][0:23], multi17 [0:24][0:23], multi18 [0:24][0:23], multi19 [0:24][0:23], multi20 [0:24][0:23], multi21 [0:24][0:23], multi22 [0:24][0:23], multi23 [0:24][0:23], multi24 [0:24][0:23];
  wire [FP_LENGTH - 1:0] sum0 [0:23][0:23], sum1 [0:23][0:23], sum2 [0:23][0:23], sum3 [0:23][0:23], sum4 [0:23][0:23], sum5 [0:23][0:23], sum6 [0:23][0:23], sum7 [0:23][0:23], sum8 [0:23][0:23], sum9 [0:23][0:23], sum10 [0:23][0:23], sum11 [0:23][0:23], sum12 [0:23][0:23], sum13 [0:23][0:23], sum14 [0:23][0:23], sum15 [0:23][0:23], sum16 [0:23][0:23], sum17 [0:23][0:23], sum18 [0:23][0:23], sum19 [0:23][0:23], sum20 [0:23][0:23], sum21 [0:23][0:23], sum22 [0:23][0:23], sum23 [0:23][0:23], sum24 [0:23][0:23];
  
//  initial begin
//    for (a = 0; a < 28; a = a + 1) begin
//        for (b = 0; b < 28; b = b + 1) begin
//            for (c = 15; c >= 0; c = c - 1) begin
//                data_array[a][b][c] = data[c + b*16 + a*28*16];
//            end
//        end
//    end
//  end
  
  genvar i0, i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21, i22, i23, m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15,m16,m17,m18,m19,m20,m21,m22,m23,m24,m25,m26,m27,m28,m29,m30,m31,m32,m33,m34,m35,m36,m37,m38,m39,m40,m41,m42,m43,m44,m45,m46,m47,m48,m49,m50,m51,m52,m53,m54,m55,m56,m57,m58,m59,m60,m61,m62,m63,m64,m65,m66,m67,m68,m69,m70,m71,m72,m73,m74,m75,m76,m77,m78,m79,m80,m81,m82,m83,m84,m85,m86,m87,m88,m89,m90,m91,m92,m93,m94,m95,m96,m97,m98,m99,m100,m101,m102,m103,m104,m105,m106,m107,m108,m109,m110,m111,m112,m113,m114,m115,m116,m117,m118,m119,m120,m121,m122,m123,m124,m125,m126,m127,m128,m129,m130,m131,m132,m133,m134,m135,m136,m137,m138,m139,m140,m141,m142,m143,m144,m145,m146,m147,m148,m149,m150,m151,m152,m153,m154,m155,m156,m157,m158,m159,m160,m161,m162,m163,m164,m165,m166,m167,m168,m169,m170,m171,m172,m173,m174,m175,m176,m177,m178,m179,m180,m181,m182,m183,m184,m185,m186,m187,m188,m189,m190,m191,m192,m193,m194,m195,m196,m197,m198,m199,m200,m201,m202,m203,m204,m205,m206,m207,m208,m209,m210,m211,m212,m213,m214,m215,m216,m217,m218,m219,m220,m221,m222,m223,m224,m225,m226,m227,m228,m229,m230,m231,m232,m233,m234,m235,m236,m237,m238,m239,m240,m241,m242,m243,m244,m245,m246,m247,m248,m249,m250,m251,m252,m253,m254,m255,m256,m257,m258,m259,m260,m261,m262,m263,m264,m265,m266,m267,m268,m269,m270,m271,m272,m273,m274,m275,m276,m277,m278,m279,m280,m281,m282,m283,m284,m285,m286,m287,m288,m289,m290,m291,m292,m293,m294,m295,m296,m297,m298,m299,m300,m301,m302,m303,m304,m305,m306,m307,m308,m309,m310,m311,m312,m313,m314,m315,m316,m317,m318,m319,m320,m321,m322,m323,m324,m325,m326,m327,m328,m329,m330,m331,m332,m333,m334,m335,m336,m337,m338,m339,m340,m341,m342,m343,m344,m345,m346,m347,m348,m349,m350,m351,m352,m353,m354,m355,m356,m357,m358,m359,m360,m361,m362,m363,m364,m365,m366,m367,m368,m369,m370,m371,m372,m373,m374,m375,m376,m377,m378,m379,m380,m381,m382,m383,m384,m385,m386,m387,m388,m389,m390,m391,m392,m393,m394,m395,m396,m397,m398,m399,m400,m401,m402,m403,m404,m405,m406,m407,m408,m409,m410,m411,m412,m413,m414,m415,m416,m417,m418,m419,m420,m421,m422,m423,m424,m425,m426,m427,m428,m429,m430,m431,m432,m433,m434,m435,m436,m437,m438,m439,m440,m441,m442,m443,m444,m445,m446,m447,m448,m449,m450,m451,m452,m453,m454,m455,m456,m457,m458,m459,m460,m461,m462,m463,m464,m465,m466,m467,m468,m469,m470,m471,m472,m473,m474,m475,m476,m477,m478,m479,m480,m481,m482,m483,m484,m485,m486,m487,m488,m489,m490,m491,m492,m493,m494,m495,m496,m497,m498,m499,m500,m501,m502,m503,m504,m505,m506,m507,m508,m509,m510,m511,m512,m513,m514,m515,m516,m517,m518,m519,m520,m521,m522,m523,m524,m525,m526,m527,m528,m529,m530,m531,m532,m533,m534,m535,m536,m537,m538,m539,m540,m541,m542,m543,m544,m545,m546,m547,m548,m549,m550,m551,m552,m553,m554,m555,m556,m557,m558,m559,m560,m561,m562,m563,m564,m565,m566,m567,m568,m569,m570,m571,m572,m573,m574,m575,m576,m577,m578,m579,m580,m581,m582,m583,m584,m585,m586,m587,m588,m589,m590,m591,m592,m593,m594,m595,m596,m597,m598,m599,m600,m601,m602,m603,m604,m605,m606,m607,m608,m609,m610,m611,m612,m613,m614,m615,m616,m617,m618,m619,m620,m621,m622,m623,m624,m625,m626,m627,m628,m629,m630,m631,m632,m633,m634,m635,m636,m637,m638,m639,m640,m641,m642,m643,m644,m645,m646,m647,m648,m649,m650,m651,m652,m653,m654,m655,m656,m657,m658,m659,m660,m661,m662,m663,m664,m665,m666,m667,m668,m669,m670,m671,m672,m673,m674,m675,m676,m677,m678,m679,m680,m681,m682,m683,m684,m685,m686,m687,m688,m689,m690,m691,m692,m693,m694,m695,m696,m697,m698,m699,m700,m701,m702,m703,m704,m705,m706,m707,m708,m709,m710,m711,m712,m713,m714,m715,m716,m717,m718,m719,m720,m721,m722,m723,m724,m725,m726,m727,m728,m729,m730,m731,m732,m733,m734,m735,m736,m737,m738,m739,m740,m741,m742,m743,m744,m745,m746,m747,m748,m749,m750,m751,m752,m753,m754,m755,m756,m757,m758,m759,m760,m761,m762,m763,m764,m765,m766,m767,m768,m769,m770,m771,m772,m773,m774,m775,m776,m777,m778,m779,m780,m781,m782,m783,n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n50,n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80,n81,n82,n83,n84,n85,n86,n87,n88,n89,n90,n91,n92,n93,n94,n95,n96,n97,n98,n99,n100,n101,n102,n103,n104,n105,n106,n107,n108,n109,n110,n111,n112,n113,n114,n115,n116,n117,n118,n119,n120,n121,n122,n123,n124,n125,n126,n127,n128,n129,n130,n131,n132,n133,n134,n135,n136,n137,n138,n139,n140,n141,n142,n143,n144,n145,n146,n147,n148,n149,n150,n151,n152,n153,n154,n155,n156,n157,n158,n159,n160,n161,n162,n163,n164,n165,n166,n167,n168,n169,n170,n171,n172,n173,n174,n175,n176,n177,n178,n179,n180,n181,n182,n183,n184,n185,n186,n187,n188,n189,n190,n191,n192,n193,n194,n195,n196,n197,n198,n199,n200,n201,n202,n203,n204,n205,n206,n207,n208,n209,n210,n211,n212,n213,n214,n215,n216,n217,n218,n219,n220,n221,n222,n223,n224,n225,n226,n227,n228,n229,n230,n231,n232,n233,n234,n235,n236,n237,n238,n239,n240,n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,n251,n252,n253,n254,n255,n256,n257,n258,n259,n260,n261,n262,n263,n264,n265,n266,n267,n268,n269,n270,n271,n272,n273,n274,n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,n330,n331,n332,n333,n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,n345,n346,n347,n348,n349,n350,n351,n352,n353,n354,n355,n356,n357,n358,n359,n360,n361,n362,n363,n364,n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,n385,n386,n387,n388,n389,n390,n391,n392,n393,n394,n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,n415,n416,n417,n418,n419,n420,n421,n422,n423,n424,n425,n426,n427,n428,n429,n430,n431,n432,n433,n434,n435,n436,n437,n438,n439,n440,n441,n442,n443,n444,n445,n446,n447,n448,n449,n450,n451,n452,n453,n454,n455,n456,n457,n458,n459,n460,n461,n462,n463,n464,n465,n466,n467,n468,n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,n479,n480,n481,n482,n483,n484,n485,n486,n487,n488,n489,n490,n491,n492,n493,n494,n495,n496,n497,n498,n499,n500,n501,n502,n503,n504,n505,n506,n507,n508,n509,n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,n559,n560,n561,n562,n563,n564,n565,n566,n567,n568,n569,n570,n571,n572,n573,n574,n575,n576,n577,n578,n579,n580,n581,n582,n583,n584,n585,n586,n587,n588,n589,n590,n591,n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,n612,n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,n623,n624,n625,n626,n627,n628,n629,n630,n631,n632,n633,n634,n635,n636,n637,n638,n639,n640,n641,n642,n643,n644,n645,n646,n647,n648,n649,n650,n651,n652,n653,n654,n655,n656,n657,n658,n659,n660,n661,n662,n663,n664,n665,n666,n667,n668,n669,n670,n671,n672,n673,n674,n675,n676,n677,n678,n679,n680,n681,n682,n683,n684,n685,n686,n687,n688,n689,n690,n691,n692,n693,n694,n695,n696,n697,n698,n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,n709,n710,n711,n712,n713,n714,n715,n716,n717,n718,n719,n720,n721,n722,n723,n724,n725,n726,n727,n728,n729,n730,n731,n732,n733,n734,n735,n736,n737,n738,n739,n740,n741,n742,n743,n744,n745,n746,n747,n748,n749,n750,n751,n752,n753,n754,n755,n756,n757,n758,n759,n760,n761,n762,n763,n764,n765,n766,n767,n768,n769,n770,n771,n772,n773,n774,n775,n776,n777,n778,n779,n780,n781,n782,n783;
  
  localparam integer a0 = 0;
    generate 
        localparam integer b0 = 0;
        for (m0 = 0; m0 < 16; m0 = m0 + 1) 
        begin: inbit0
            assign data_11[m0 + b0*16 + a0*28*16] = data_11_array[a0][b0][m0];
        end
    endgenerate
    generate 
        localparam integer b1 = 1;
        for (m1 = 0; m1 < 16; m1 = m1 + 1) 
        begin: inbit1
            assign data_11[m1 + b1*16 + a0*28*16] = data_11_array[a0][b1][m1];
        end
    endgenerate
    generate 
        localparam integer b2 = 2;
        for (m2 = 0; m2 < 16; m2 = m2 + 1) 
        begin: inbit2
            assign data_11[m2 + b2*16 + a0*28*16] = data_11_array[a0][b2][m2];
        end
    endgenerate
    generate 
        localparam integer b3 = 3;
        for (m3 = 0; m3 < 16; m3 = m3 + 1) 
        begin: inbit3
            assign data_11[m3 + b3*16 + a0*28*16] = data_11_array[a0][b3][m3];
        end
    endgenerate
    generate 
        localparam integer b4 = 4;
        for (m4 = 0; m4 < 16; m4 = m4 + 1) 
        begin: inbit4
            assign data_11[m4 + b4*16 + a0*28*16] = data_11_array[a0][b4][m4];
        end
    endgenerate
    generate 
        localparam integer b5 = 5;
        for (m5 = 0; m5 < 16; m5 = m5 + 1) 
        begin: inbit5
            assign data_11[m5 + b5*16 + a0*28*16] = data_11_array[a0][b5][m5];
        end
    endgenerate
    generate 
        localparam integer b6 = 6;
        for (m6 = 0; m6 < 16; m6 = m6 + 1) 
        begin: inbit6
            assign data_11[m6 + b6*16 + a0*28*16] = data_11_array[a0][b6][m6];
        end
    endgenerate
    generate 
        localparam integer b7 = 7;
        for (m7 = 0; m7 < 16; m7 = m7 + 1) 
        begin: inbit7
            assign data_11[m7 + b7*16 + a0*28*16] = data_11_array[a0][b7][m7];
        end
    endgenerate
    generate 
        localparam integer b8 = 8;
        for (m8 = 0; m8 < 16; m8 = m8 + 1) 
        begin: inbit8
            assign data_11[m8 + b8*16 + a0*28*16] = data_11_array[a0][b8][m8];
        end
    endgenerate
    generate 
        localparam integer b9 = 9;
        for (m9 = 0; m9 < 16; m9 = m9 + 1) 
        begin: inbit9
            assign data_11[m9 + b9*16 + a0*28*16] = data_11_array[a0][b9][m9];
        end
    endgenerate
    generate 
        localparam integer b10 = 10;
        for (m10 = 0; m10 < 16; m10 = m10 + 1) 
        begin: inbit10
            assign data_11[m10 + b10*16 + a0*28*16] = data_11_array[a0][b10][m10];
        end
    endgenerate
    generate 
        localparam integer b11 = 11;
        for (m11 = 0; m11 < 16; m11 = m11 + 1) 
        begin: inbit11
            assign data_11[m11 + b11*16 + a0*28*16] = data_11_array[a0][b11][m11];
        end
    endgenerate
    generate 
        localparam integer b12 = 12;
        for (m12 = 0; m12 < 16; m12 = m12 + 1) 
        begin: inbit12
            assign data_11[m12 + b12*16 + a0*28*16] = data_11_array[a0][b12][m12];
        end
    endgenerate
    generate 
        localparam integer b13 = 13;
        for (m13 = 0; m13 < 16; m13 = m13 + 1) 
        begin: inbit13
            assign data_11[m13 + b13*16 + a0*28*16] = data_11_array[a0][b13][m13];
        end
    endgenerate
    generate 
        localparam integer b14 = 14;
        for (m14 = 0; m14 < 16; m14 = m14 + 1) 
        begin: inbit14
            assign data_11[m14 + b14*16 + a0*28*16] = data_11_array[a0][b14][m14];
        end
    endgenerate
    generate 
        localparam integer b15 = 15;
        for (m15 = 0; m15 < 16; m15 = m15 + 1) 
        begin: inbit15
            assign data_11[m15 + b15*16 + a0*28*16] = data_11_array[a0][b15][m15];
        end
    endgenerate
    generate 
        localparam integer b16 = 16;
        for (m16 = 0; m16 < 16; m16 = m16 + 1) 
        begin: inbit16
            assign data_11[m16 + b16*16 + a0*28*16] = data_11_array[a0][b16][m16];
        end
    endgenerate
    generate 
        localparam integer b17 = 17;
        for (m17 = 0; m17 < 16; m17 = m17 + 1) 
        begin: inbit17
            assign data_11[m17 + b17*16 + a0*28*16] = data_11_array[a0][b17][m17];
        end
    endgenerate
    generate 
        localparam integer b18 = 18;
        for (m18 = 0; m18 < 16; m18 = m18 + 1) 
        begin: inbit18
            assign data_11[m18 + b18*16 + a0*28*16] = data_11_array[a0][b18][m18];
        end
    endgenerate
    generate 
        localparam integer b19 = 19;
        for (m19 = 0; m19 < 16; m19 = m19 + 1) 
        begin: inbit19
            assign data_11[m19 + b19*16 + a0*28*16] = data_11_array[a0][b19][m19];
        end
    endgenerate
    generate 
        localparam integer b20 = 20;
        for (m20 = 0; m20 < 16; m20 = m20 + 1) 
        begin: inbit20
            assign data_11[m20 + b20*16 + a0*28*16] = data_11_array[a0][b20][m20];
        end
    endgenerate
    generate 
        localparam integer b21 = 21;
        for (m21 = 0; m21 < 16; m21 = m21 + 1) 
        begin: inbit21
            assign data_11[m21 + b21*16 + a0*28*16] = data_11_array[a0][b21][m21];
        end
    endgenerate
    generate 
        localparam integer b22 = 22;
        for (m22 = 0; m22 < 16; m22 = m22 + 1) 
        begin: inbit22
            assign data_11[m22 + b22*16 + a0*28*16] = data_11_array[a0][b22][m22];
        end
    endgenerate
    generate 
        localparam integer b23 = 23;
        for (m23 = 0; m23 < 16; m23 = m23 + 1) 
        begin: inbit23
            assign data_11[m23 + b23*16 + a0*28*16] = data_11_array[a0][b23][m23];
        end
    endgenerate
    generate 
        localparam integer b24 = 24;
        for (m24 = 0; m24 < 16; m24 = m24 + 1) 
        begin: inbit24
            assign data_11[m24 + b24*16 + a0*28*16] = data_11_array[a0][b24][m24];
        end
    endgenerate
    generate 
        localparam integer b25 = 25;
        for (m25 = 0; m25 < 16; m25 = m25 + 1) 
        begin: inbit25
            assign data_11[m25 + b25*16 + a0*28*16] = data_11_array[a0][b25][m25];
        end
    endgenerate
    generate 
        localparam integer b26 = 26;
        for (m26 = 0; m26 < 16; m26 = m26 + 1) 
        begin: inbit26
            assign data_11[m26 + b26*16 + a0*28*16] = data_11_array[a0][b26][m26];
        end
    endgenerate
    generate 
        localparam integer b27 = 27;
        for (m27 = 0; m27 < 16; m27 = m27 + 1) 
        begin: inbit27
            assign data_11[m27 + b27*16 + a0*28*16] = data_11_array[a0][b27][m27];
        end
    endgenerate
    localparam integer a1 = 1;
    generate 
        localparam integer b28 = 0;
        for (m28 = 0; m28 < 16; m28 = m28 + 1) 
        begin: inbit28
            assign data_11[m28 + b28*16 + a1*28*16] = data_11_array[a1][b28][m28];
        end
    endgenerate
    generate 
        localparam integer b29 = 1;
        for (m29 = 0; m29 < 16; m29 = m29 + 1) 
        begin: inbit29
            assign data_11[m29 + b29*16 + a1*28*16] = data_11_array[a1][b29][m29];
        end
    endgenerate
    generate 
        localparam integer b30 = 2;
        for (m30 = 0; m30 < 16; m30 = m30 + 1) 
        begin: inbit30
            assign data_11[m30 + b30*16 + a1*28*16] = data_11_array[a1][b30][m30];
        end
    endgenerate
    generate 
        localparam integer b31 = 3;
        for (m31 = 0; m31 < 16; m31 = m31 + 1) 
        begin: inbit31
            assign data_11[m31 + b31*16 + a1*28*16] = data_11_array[a1][b31][m31];
        end
    endgenerate
    generate 
        localparam integer b32 = 4;
        for (m32 = 0; m32 < 16; m32 = m32 + 1) 
        begin: inbit32
            assign data_11[m32 + b32*16 + a1*28*16] = data_11_array[a1][b32][m32];
        end
    endgenerate
    generate 
        localparam integer b33 = 5;
        for (m33 = 0; m33 < 16; m33 = m33 + 1) 
        begin: inbit33
            assign data_11[m33 + b33*16 + a1*28*16] = data_11_array[a1][b33][m33];
        end
    endgenerate
    generate 
        localparam integer b34 = 6;
        for (m34 = 0; m34 < 16; m34 = m34 + 1) 
        begin: inbit34
            assign data_11[m34 + b34*16 + a1*28*16] = data_11_array[a1][b34][m34];
        end
    endgenerate
    generate 
        localparam integer b35 = 7;
        for (m35 = 0; m35 < 16; m35 = m35 + 1) 
        begin: inbit35
            assign data_11[m35 + b35*16 + a1*28*16] = data_11_array[a1][b35][m35];
        end
    endgenerate
    generate 
        localparam integer b36 = 8;
        for (m36 = 0; m36 < 16; m36 = m36 + 1) 
        begin: inbit36
            assign data_11[m36 + b36*16 + a1*28*16] = data_11_array[a1][b36][m36];
        end
    endgenerate
    generate 
        localparam integer b37 = 9;
        for (m37 = 0; m37 < 16; m37 = m37 + 1) 
        begin: inbit37
            assign data_11[m37 + b37*16 + a1*28*16] = data_11_array[a1][b37][m37];
        end
    endgenerate
    generate 
        localparam integer b38 = 10;
        for (m38 = 0; m38 < 16; m38 = m38 + 1) 
        begin: inbit38
            assign data_11[m38 + b38*16 + a1*28*16] = data_11_array[a1][b38][m38];
        end
    endgenerate
    generate 
        localparam integer b39 = 11;
        for (m39 = 0; m39 < 16; m39 = m39 + 1) 
        begin: inbit39
            assign data_11[m39 + b39*16 + a1*28*16] = data_11_array[a1][b39][m39];
        end
    endgenerate
    generate 
        localparam integer b40 = 12;
        for (m40 = 0; m40 < 16; m40 = m40 + 1) 
        begin: inbit40
            assign data_11[m40 + b40*16 + a1*28*16] = data_11_array[a1][b40][m40];
        end
    endgenerate
    generate 
        localparam integer b41 = 13;
        for (m41 = 0; m41 < 16; m41 = m41 + 1) 
        begin: inbit41
            assign data_11[m41 + b41*16 + a1*28*16] = data_11_array[a1][b41][m41];
        end
    endgenerate
    generate 
        localparam integer b42 = 14;
        for (m42 = 0; m42 < 16; m42 = m42 + 1) 
        begin: inbit42
            assign data_11[m42 + b42*16 + a1*28*16] = data_11_array[a1][b42][m42];
        end
    endgenerate
    generate 
        localparam integer b43 = 15;
        for (m43 = 0; m43 < 16; m43 = m43 + 1) 
        begin: inbit43
            assign data_11[m43 + b43*16 + a1*28*16] = data_11_array[a1][b43][m43];
        end
    endgenerate
    generate 
        localparam integer b44 = 16;
        for (m44 = 0; m44 < 16; m44 = m44 + 1) 
        begin: inbit44
            assign data_11[m44 + b44*16 + a1*28*16] = data_11_array[a1][b44][m44];
        end
    endgenerate
    generate 
        localparam integer b45 = 17;
        for (m45 = 0; m45 < 16; m45 = m45 + 1) 
        begin: inbit45
            assign data_11[m45 + b45*16 + a1*28*16] = data_11_array[a1][b45][m45];
        end
    endgenerate
    generate 
        localparam integer b46 = 18;
        for (m46 = 0; m46 < 16; m46 = m46 + 1) 
        begin: inbit46
            assign data_11[m46 + b46*16 + a1*28*16] = data_11_array[a1][b46][m46];
        end
    endgenerate
    generate 
        localparam integer b47 = 19;
        for (m47 = 0; m47 < 16; m47 = m47 + 1) 
        begin: inbit47
            assign data_11[m47 + b47*16 + a1*28*16] = data_11_array[a1][b47][m47];
        end
    endgenerate
    generate 
        localparam integer b48 = 20;
        for (m48 = 0; m48 < 16; m48 = m48 + 1) 
        begin: inbit48
            assign data_11[m48 + b48*16 + a1*28*16] = data_11_array[a1][b48][m48];
        end
    endgenerate
    generate 
        localparam integer b49 = 21;
        for (m49 = 0; m49 < 16; m49 = m49 + 1) 
        begin: inbit49
            assign data_11[m49 + b49*16 + a1*28*16] = data_11_array[a1][b49][m49];
        end
    endgenerate
    generate 
        localparam integer b50 = 22;
        for (m50 = 0; m50 < 16; m50 = m50 + 1) 
        begin: inbit50
            assign data_11[m50 + b50*16 + a1*28*16] = data_11_array[a1][b50][m50];
        end
    endgenerate
    generate 
        localparam integer b51 = 23;
        for (m51 = 0; m51 < 16; m51 = m51 + 1) 
        begin: inbit51
            assign data_11[m51 + b51*16 + a1*28*16] = data_11_array[a1][b51][m51];
        end
    endgenerate
    generate 
        localparam integer b52 = 24;
        for (m52 = 0; m52 < 16; m52 = m52 + 1) 
        begin: inbit52
            assign data_11[m52 + b52*16 + a1*28*16] = data_11_array[a1][b52][m52];
        end
    endgenerate
    generate 
        localparam integer b53 = 25;
        for (m53 = 0; m53 < 16; m53 = m53 + 1) 
        begin: inbit53
            assign data_11[m53 + b53*16 + a1*28*16] = data_11_array[a1][b53][m53];
        end
    endgenerate
    generate 
        localparam integer b54 = 26;
        for (m54 = 0; m54 < 16; m54 = m54 + 1) 
        begin: inbit54
            assign data_11[m54 + b54*16 + a1*28*16] = data_11_array[a1][b54][m54];
        end
    endgenerate
    generate 
        localparam integer b55 = 27;
        for (m55 = 0; m55 < 16; m55 = m55 + 1) 
        begin: inbit55
            assign data_11[m55 + b55*16 + a1*28*16] = data_11_array[a1][b55][m55];
        end
    endgenerate
    localparam integer a2 = 2;
    generate 
        localparam integer b56 = 0;
        for (m56 = 0; m56 < 16; m56 = m56 + 1) 
        begin: inbit56
            assign data_11[m56 + b56*16 + a2*28*16] = data_11_array[a2][b56][m56];
        end
    endgenerate
    generate 
        localparam integer b57 = 1;
        for (m57 = 0; m57 < 16; m57 = m57 + 1) 
        begin: inbit57
            assign data_11[m57 + b57*16 + a2*28*16] = data_11_array[a2][b57][m57];
        end
    endgenerate
    generate 
        localparam integer b58 = 2;
        for (m58 = 0; m58 < 16; m58 = m58 + 1) 
        begin: inbit58
            assign data_11[m58 + b58*16 + a2*28*16] = data_11_array[a2][b58][m58];
        end
    endgenerate
    generate 
        localparam integer b59 = 3;
        for (m59 = 0; m59 < 16; m59 = m59 + 1) 
        begin: inbit59
            assign data_11[m59 + b59*16 + a2*28*16] = data_11_array[a2][b59][m59];
        end
    endgenerate
    generate 
        localparam integer b60 = 4;
        for (m60 = 0; m60 < 16; m60 = m60 + 1) 
        begin: inbit60
            assign data_11[m60 + b60*16 + a2*28*16] = data_11_array[a2][b60][m60];
        end
    endgenerate
    generate 
        localparam integer b61 = 5;
        for (m61 = 0; m61 < 16; m61 = m61 + 1) 
        begin: inbit61
            assign data_11[m61 + b61*16 + a2*28*16] = data_11_array[a2][b61][m61];
        end
    endgenerate
    generate 
        localparam integer b62 = 6;
        for (m62 = 0; m62 < 16; m62 = m62 + 1) 
        begin: inbit62
            assign data_11[m62 + b62*16 + a2*28*16] = data_11_array[a2][b62][m62];
        end
    endgenerate
    generate 
        localparam integer b63 = 7;
        for (m63 = 0; m63 < 16; m63 = m63 + 1) 
        begin: inbit63
            assign data_11[m63 + b63*16 + a2*28*16] = data_11_array[a2][b63][m63];
        end
    endgenerate
    generate 
        localparam integer b64 = 8;
        for (m64 = 0; m64 < 16; m64 = m64 + 1) 
        begin: inbit64
            assign data_11[m64 + b64*16 + a2*28*16] = data_11_array[a2][b64][m64];
        end
    endgenerate
    generate 
        localparam integer b65 = 9;
        for (m65 = 0; m65 < 16; m65 = m65 + 1) 
        begin: inbit65
            assign data_11[m65 + b65*16 + a2*28*16] = data_11_array[a2][b65][m65];
        end
    endgenerate
    generate 
        localparam integer b66 = 10;
        for (m66 = 0; m66 < 16; m66 = m66 + 1) 
        begin: inbit66
            assign data_11[m66 + b66*16 + a2*28*16] = data_11_array[a2][b66][m66];
        end
    endgenerate
    generate 
        localparam integer b67 = 11;
        for (m67 = 0; m67 < 16; m67 = m67 + 1) 
        begin: inbit67
            assign data_11[m67 + b67*16 + a2*28*16] = data_11_array[a2][b67][m67];
        end
    endgenerate
    generate 
        localparam integer b68 = 12;
        for (m68 = 0; m68 < 16; m68 = m68 + 1) 
        begin: inbit68
            assign data_11[m68 + b68*16 + a2*28*16] = data_11_array[a2][b68][m68];
        end
    endgenerate
    generate 
        localparam integer b69 = 13;
        for (m69 = 0; m69 < 16; m69 = m69 + 1) 
        begin: inbit69
            assign data_11[m69 + b69*16 + a2*28*16] = data_11_array[a2][b69][m69];
        end
    endgenerate
    generate 
        localparam integer b70 = 14;
        for (m70 = 0; m70 < 16; m70 = m70 + 1) 
        begin: inbit70
            assign data_11[m70 + b70*16 + a2*28*16] = data_11_array[a2][b70][m70];
        end
    endgenerate
    generate 
        localparam integer b71 = 15;
        for (m71 = 0; m71 < 16; m71 = m71 + 1) 
        begin: inbit71
            assign data_11[m71 + b71*16 + a2*28*16] = data_11_array[a2][b71][m71];
        end
    endgenerate
    generate 
        localparam integer b72 = 16;
        for (m72 = 0; m72 < 16; m72 = m72 + 1) 
        begin: inbit72
            assign data_11[m72 + b72*16 + a2*28*16] = data_11_array[a2][b72][m72];
        end
    endgenerate
    generate 
        localparam integer b73 = 17;
        for (m73 = 0; m73 < 16; m73 = m73 + 1) 
        begin: inbit73
            assign data_11[m73 + b73*16 + a2*28*16] = data_11_array[a2][b73][m73];
        end
    endgenerate
    generate 
        localparam integer b74 = 18;
        for (m74 = 0; m74 < 16; m74 = m74 + 1) 
        begin: inbit74
            assign data_11[m74 + b74*16 + a2*28*16] = data_11_array[a2][b74][m74];
        end
    endgenerate
    generate 
        localparam integer b75 = 19;
        for (m75 = 0; m75 < 16; m75 = m75 + 1) 
        begin: inbit75
            assign data_11[m75 + b75*16 + a2*28*16] = data_11_array[a2][b75][m75];
        end
    endgenerate
    generate 
        localparam integer b76 = 20;
        for (m76 = 0; m76 < 16; m76 = m76 + 1) 
        begin: inbit76
            assign data_11[m76 + b76*16 + a2*28*16] = data_11_array[a2][b76][m76];
        end
    endgenerate
    generate 
        localparam integer b77 = 21;
        for (m77 = 0; m77 < 16; m77 = m77 + 1) 
        begin: inbit77
            assign data_11[m77 + b77*16 + a2*28*16] = data_11_array[a2][b77][m77];
        end
    endgenerate
    generate 
        localparam integer b78 = 22;
        for (m78 = 0; m78 < 16; m78 = m78 + 1) 
        begin: inbit78
            assign data_11[m78 + b78*16 + a2*28*16] = data_11_array[a2][b78][m78];
        end
    endgenerate
    generate 
        localparam integer b79 = 23;
        for (m79 = 0; m79 < 16; m79 = m79 + 1) 
        begin: inbit79
            assign data_11[m79 + b79*16 + a2*28*16] = data_11_array[a2][b79][m79];
        end
    endgenerate
    generate 
        localparam integer b80 = 24;
        for (m80 = 0; m80 < 16; m80 = m80 + 1) 
        begin: inbit80
            assign data_11[m80 + b80*16 + a2*28*16] = data_11_array[a2][b80][m80];
        end
    endgenerate
    generate 
        localparam integer b81 = 25;
        for (m81 = 0; m81 < 16; m81 = m81 + 1) 
        begin: inbit81
            assign data_11[m81 + b81*16 + a2*28*16] = data_11_array[a2][b81][m81];
        end
    endgenerate
    generate 
        localparam integer b82 = 26;
        for (m82 = 0; m82 < 16; m82 = m82 + 1) 
        begin: inbit82
            assign data_11[m82 + b82*16 + a2*28*16] = data_11_array[a2][b82][m82];
        end
    endgenerate
    generate 
        localparam integer b83 = 27;
        for (m83 = 0; m83 < 16; m83 = m83 + 1) 
        begin: inbit83
            assign data_11[m83 + b83*16 + a2*28*16] = data_11_array[a2][b83][m83];
        end
    endgenerate
    localparam integer a3 = 3;
    generate 
        localparam integer b84 = 0;
        for (m84 = 0; m84 < 16; m84 = m84 + 1) 
        begin: inbit84
            assign data_11[m84 + b84*16 + a3*28*16] = data_11_array[a3][b84][m84];
        end
    endgenerate
    generate 
        localparam integer b85 = 1;
        for (m85 = 0; m85 < 16; m85 = m85 + 1) 
        begin: inbit85
            assign data_11[m85 + b85*16 + a3*28*16] = data_11_array[a3][b85][m85];
        end
    endgenerate
    generate 
        localparam integer b86 = 2;
        for (m86 = 0; m86 < 16; m86 = m86 + 1) 
        begin: inbit86
            assign data_11[m86 + b86*16 + a3*28*16] = data_11_array[a3][b86][m86];
        end
    endgenerate
    generate 
        localparam integer b87 = 3;
        for (m87 = 0; m87 < 16; m87 = m87 + 1) 
        begin: inbit87
            assign data_11[m87 + b87*16 + a3*28*16] = data_11_array[a3][b87][m87];
        end
    endgenerate
    generate 
        localparam integer b88 = 4;
        for (m88 = 0; m88 < 16; m88 = m88 + 1) 
        begin: inbit88
            assign data_11[m88 + b88*16 + a3*28*16] = data_11_array[a3][b88][m88];
        end
    endgenerate
    generate 
        localparam integer b89 = 5;
        for (m89 = 0; m89 < 16; m89 = m89 + 1) 
        begin: inbit89
            assign data_11[m89 + b89*16 + a3*28*16] = data_11_array[a3][b89][m89];
        end
    endgenerate
    generate 
        localparam integer b90 = 6;
        for (m90 = 0; m90 < 16; m90 = m90 + 1) 
        begin: inbit90
            assign data_11[m90 + b90*16 + a3*28*16] = data_11_array[a3][b90][m90];
        end
    endgenerate
    generate 
        localparam integer b91 = 7;
        for (m91 = 0; m91 < 16; m91 = m91 + 1) 
        begin: inbit91
            assign data_11[m91 + b91*16 + a3*28*16] = data_11_array[a3][b91][m91];
        end
    endgenerate
    generate 
        localparam integer b92 = 8;
        for (m92 = 0; m92 < 16; m92 = m92 + 1) 
        begin: inbit92
            assign data_11[m92 + b92*16 + a3*28*16] = data_11_array[a3][b92][m92];
        end
    endgenerate
    generate 
        localparam integer b93 = 9;
        for (m93 = 0; m93 < 16; m93 = m93 + 1) 
        begin: inbit93
            assign data_11[m93 + b93*16 + a3*28*16] = data_11_array[a3][b93][m93];
        end
    endgenerate
    generate 
        localparam integer b94 = 10;
        for (m94 = 0; m94 < 16; m94 = m94 + 1) 
        begin: inbit94
            assign data_11[m94 + b94*16 + a3*28*16] = data_11_array[a3][b94][m94];
        end
    endgenerate
    generate 
        localparam integer b95 = 11;
        for (m95 = 0; m95 < 16; m95 = m95 + 1) 
        begin: inbit95
            assign data_11[m95 + b95*16 + a3*28*16] = data_11_array[a3][b95][m95];
        end
    endgenerate
    generate 
        localparam integer b96 = 12;
        for (m96 = 0; m96 < 16; m96 = m96 + 1) 
        begin: inbit96
            assign data_11[m96 + b96*16 + a3*28*16] = data_11_array[a3][b96][m96];
        end
    endgenerate
    generate 
        localparam integer b97 = 13;
        for (m97 = 0; m97 < 16; m97 = m97 + 1) 
        begin: inbit97
            assign data_11[m97 + b97*16 + a3*28*16] = data_11_array[a3][b97][m97];
        end
    endgenerate
    generate 
        localparam integer b98 = 14;
        for (m98 = 0; m98 < 16; m98 = m98 + 1) 
        begin: inbit98
            assign data_11[m98 + b98*16 + a3*28*16] = data_11_array[a3][b98][m98];
        end
    endgenerate
    generate 
        localparam integer b99 = 15;
        for (m99 = 0; m99 < 16; m99 = m99 + 1) 
        begin: inbit99
            assign data_11[m99 + b99*16 + a3*28*16] = data_11_array[a3][b99][m99];
        end
    endgenerate
    generate 
        localparam integer b100 = 16;
        for (m100 = 0; m100 < 16; m100 = m100 + 1) 
        begin: inbit100
            assign data_11[m100 + b100*16 + a3*28*16] = data_11_array[a3][b100][m100];
        end
    endgenerate
    generate 
        localparam integer b101 = 17;
        for (m101 = 0; m101 < 16; m101 = m101 + 1) 
        begin: inbit101
            assign data_11[m101 + b101*16 + a3*28*16] = data_11_array[a3][b101][m101];
        end
    endgenerate
    generate 
        localparam integer b102 = 18;
        for (m102 = 0; m102 < 16; m102 = m102 + 1) 
        begin: inbit102
            assign data_11[m102 + b102*16 + a3*28*16] = data_11_array[a3][b102][m102];
        end
    endgenerate
    generate 
        localparam integer b103 = 19;
        for (m103 = 0; m103 < 16; m103 = m103 + 1) 
        begin: inbit103
            assign data_11[m103 + b103*16 + a3*28*16] = data_11_array[a3][b103][m103];
        end
    endgenerate
    generate 
        localparam integer b104 = 20;
        for (m104 = 0; m104 < 16; m104 = m104 + 1) 
        begin: inbit104
            assign data_11[m104 + b104*16 + a3*28*16] = data_11_array[a3][b104][m104];
        end
    endgenerate
    generate 
        localparam integer b105 = 21;
        for (m105 = 0; m105 < 16; m105 = m105 + 1) 
        begin: inbit105
            assign data_11[m105 + b105*16 + a3*28*16] = data_11_array[a3][b105][m105];
        end
    endgenerate
    generate 
        localparam integer b106 = 22;
        for (m106 = 0; m106 < 16; m106 = m106 + 1) 
        begin: inbit106
            assign data_11[m106 + b106*16 + a3*28*16] = data_11_array[a3][b106][m106];
        end
    endgenerate
    generate 
        localparam integer b107 = 23;
        for (m107 = 0; m107 < 16; m107 = m107 + 1) 
        begin: inbit107
            assign data_11[m107 + b107*16 + a3*28*16] = data_11_array[a3][b107][m107];
        end
    endgenerate
    generate 
        localparam integer b108 = 24;
        for (m108 = 0; m108 < 16; m108 = m108 + 1) 
        begin: inbit108
            assign data_11[m108 + b108*16 + a3*28*16] = data_11_array[a3][b108][m108];
        end
    endgenerate
    generate 
        localparam integer b109 = 25;
        for (m109 = 0; m109 < 16; m109 = m109 + 1) 
        begin: inbit109
            assign data_11[m109 + b109*16 + a3*28*16] = data_11_array[a3][b109][m109];
        end
    endgenerate
    generate 
        localparam integer b110 = 26;
        for (m110 = 0; m110 < 16; m110 = m110 + 1) 
        begin: inbit110
            assign data_11[m110 + b110*16 + a3*28*16] = data_11_array[a3][b110][m110];
        end
    endgenerate
    generate 
        localparam integer b111 = 27;
        for (m111 = 0; m111 < 16; m111 = m111 + 1) 
        begin: inbit111
            assign data_11[m111 + b111*16 + a3*28*16] = data_11_array[a3][b111][m111];
        end
    endgenerate
    localparam integer a4 = 4;
    generate 
        localparam integer b112 = 0;
        for (m112 = 0; m112 < 16; m112 = m112 + 1) 
        begin: inbit112
            assign data_11[m112 + b112*16 + a4*28*16] = data_11_array[a4][b112][m112];
        end
    endgenerate
    generate 
        localparam integer b113 = 1;
        for (m113 = 0; m113 < 16; m113 = m113 + 1) 
        begin: inbit113
            assign data_11[m113 + b113*16 + a4*28*16] = data_11_array[a4][b113][m113];
        end
    endgenerate
    generate 
        localparam integer b114 = 2;
        for (m114 = 0; m114 < 16; m114 = m114 + 1) 
        begin: inbit114
            assign data_11[m114 + b114*16 + a4*28*16] = data_11_array[a4][b114][m114];
        end
    endgenerate
    generate 
        localparam integer b115 = 3;
        for (m115 = 0; m115 < 16; m115 = m115 + 1) 
        begin: inbit115
            assign data_11[m115 + b115*16 + a4*28*16] = data_11_array[a4][b115][m115];
        end
    endgenerate
    generate 
        localparam integer b116 = 4;
        for (m116 = 0; m116 < 16; m116 = m116 + 1) 
        begin: inbit116
            assign data_11[m116 + b116*16 + a4*28*16] = data_11_array[a4][b116][m116];
        end
    endgenerate
    generate 
        localparam integer b117 = 5;
        for (m117 = 0; m117 < 16; m117 = m117 + 1) 
        begin: inbit117
            assign data_11[m117 + b117*16 + a4*28*16] = data_11_array[a4][b117][m117];
        end
    endgenerate
    generate 
        localparam integer b118 = 6;
        for (m118 = 0; m118 < 16; m118 = m118 + 1) 
        begin: inbit118
            assign data_11[m118 + b118*16 + a4*28*16] = data_11_array[a4][b118][m118];
        end
    endgenerate
    generate 
        localparam integer b119 = 7;
        for (m119 = 0; m119 < 16; m119 = m119 + 1) 
        begin: inbit119
            assign data_11[m119 + b119*16 + a4*28*16] = data_11_array[a4][b119][m119];
        end
    endgenerate
    generate 
        localparam integer b120 = 8;
        for (m120 = 0; m120 < 16; m120 = m120 + 1) 
        begin: inbit120
            assign data_11[m120 + b120*16 + a4*28*16] = data_11_array[a4][b120][m120];
        end
    endgenerate
    generate 
        localparam integer b121 = 9;
        for (m121 = 0; m121 < 16; m121 = m121 + 1) 
        begin: inbit121
            assign data_11[m121 + b121*16 + a4*28*16] = data_11_array[a4][b121][m121];
        end
    endgenerate
    generate 
        localparam integer b122 = 10;
        for (m122 = 0; m122 < 16; m122 = m122 + 1) 
        begin: inbit122
            assign data_11[m122 + b122*16 + a4*28*16] = data_11_array[a4][b122][m122];
        end
    endgenerate
    generate 
        localparam integer b123 = 11;
        for (m123 = 0; m123 < 16; m123 = m123 + 1) 
        begin: inbit123
            assign data_11[m123 + b123*16 + a4*28*16] = data_11_array[a4][b123][m123];
        end
    endgenerate
    generate 
        localparam integer b124 = 12;
        for (m124 = 0; m124 < 16; m124 = m124 + 1) 
        begin: inbit124
            assign data_11[m124 + b124*16 + a4*28*16] = data_11_array[a4][b124][m124];
        end
    endgenerate
    generate 
        localparam integer b125 = 13;
        for (m125 = 0; m125 < 16; m125 = m125 + 1) 
        begin: inbit125
            assign data_11[m125 + b125*16 + a4*28*16] = data_11_array[a4][b125][m125];
        end
    endgenerate
    generate 
        localparam integer b126 = 14;
        for (m126 = 0; m126 < 16; m126 = m126 + 1) 
        begin: inbit126
            assign data_11[m126 + b126*16 + a4*28*16] = data_11_array[a4][b126][m126];
        end
    endgenerate
    generate 
        localparam integer b127 = 15;
        for (m127 = 0; m127 < 16; m127 = m127 + 1) 
        begin: inbit127
            assign data_11[m127 + b127*16 + a4*28*16] = data_11_array[a4][b127][m127];
        end
    endgenerate
    generate 
        localparam integer b128 = 16;
        for (m128 = 0; m128 < 16; m128 = m128 + 1) 
        begin: inbit128
            assign data_11[m128 + b128*16 + a4*28*16] = data_11_array[a4][b128][m128];
        end
    endgenerate
    generate 
        localparam integer b129 = 17;
        for (m129 = 0; m129 < 16; m129 = m129 + 1) 
        begin: inbit129
            assign data_11[m129 + b129*16 + a4*28*16] = data_11_array[a4][b129][m129];
        end
    endgenerate
    generate 
        localparam integer b130 = 18;
        for (m130 = 0; m130 < 16; m130 = m130 + 1) 
        begin: inbit130
            assign data_11[m130 + b130*16 + a4*28*16] = data_11_array[a4][b130][m130];
        end
    endgenerate
    generate 
        localparam integer b131 = 19;
        for (m131 = 0; m131 < 16; m131 = m131 + 1) 
        begin: inbit131
            assign data_11[m131 + b131*16 + a4*28*16] = data_11_array[a4][b131][m131];
        end
    endgenerate
    generate 
        localparam integer b132 = 20;
        for (m132 = 0; m132 < 16; m132 = m132 + 1) 
        begin: inbit132
            assign data_11[m132 + b132*16 + a4*28*16] = data_11_array[a4][b132][m132];
        end
    endgenerate
    generate 
        localparam integer b133 = 21;
        for (m133 = 0; m133 < 16; m133 = m133 + 1) 
        begin: inbit133
            assign data_11[m133 + b133*16 + a4*28*16] = data_11_array[a4][b133][m133];
        end
    endgenerate
    generate 
        localparam integer b134 = 22;
        for (m134 = 0; m134 < 16; m134 = m134 + 1) 
        begin: inbit134
            assign data_11[m134 + b134*16 + a4*28*16] = data_11_array[a4][b134][m134];
        end
    endgenerate
    generate 
        localparam integer b135 = 23;
        for (m135 = 0; m135 < 16; m135 = m135 + 1) 
        begin: inbit135
            assign data_11[m135 + b135*16 + a4*28*16] = data_11_array[a4][b135][m135];
        end
    endgenerate
    generate 
        localparam integer b136 = 24;
        for (m136 = 0; m136 < 16; m136 = m136 + 1) 
        begin: inbit136
            assign data_11[m136 + b136*16 + a4*28*16] = data_11_array[a4][b136][m136];
        end
    endgenerate
    generate 
        localparam integer b137 = 25;
        for (m137 = 0; m137 < 16; m137 = m137 + 1) 
        begin: inbit137
            assign data_11[m137 + b137*16 + a4*28*16] = data_11_array[a4][b137][m137];
        end
    endgenerate
    generate 
        localparam integer b138 = 26;
        for (m138 = 0; m138 < 16; m138 = m138 + 1) 
        begin: inbit138
            assign data_11[m138 + b138*16 + a4*28*16] = data_11_array[a4][b138][m138];
        end
    endgenerate
    generate 
        localparam integer b139 = 27;
        for (m139 = 0; m139 < 16; m139 = m139 + 1) 
        begin: inbit139
            assign data_11[m139 + b139*16 + a4*28*16] = data_11_array[a4][b139][m139];
        end
    endgenerate
    localparam integer a5 = 5;
    generate 
        localparam integer b140 = 0;
        for (m140 = 0; m140 < 16; m140 = m140 + 1) 
        begin: inbit140
            assign data_11[m140 + b140*16 + a5*28*16] = data_11_array[a5][b140][m140];
        end
    endgenerate
    generate 
        localparam integer b141 = 1;
        for (m141 = 0; m141 < 16; m141 = m141 + 1) 
        begin: inbit141
            assign data_11[m141 + b141*16 + a5*28*16] = data_11_array[a5][b141][m141];
        end
    endgenerate
    generate 
        localparam integer b142 = 2;
        for (m142 = 0; m142 < 16; m142 = m142 + 1) 
        begin: inbit142
            assign data_11[m142 + b142*16 + a5*28*16] = data_11_array[a5][b142][m142];
        end
    endgenerate
    generate 
        localparam integer b143 = 3;
        for (m143 = 0; m143 < 16; m143 = m143 + 1) 
        begin: inbit143
            assign data_11[m143 + b143*16 + a5*28*16] = data_11_array[a5][b143][m143];
        end
    endgenerate
    generate 
        localparam integer b144 = 4;
        for (m144 = 0; m144 < 16; m144 = m144 + 1) 
        begin: inbit144
            assign data_11[m144 + b144*16 + a5*28*16] = data_11_array[a5][b144][m144];
        end
    endgenerate
    generate 
        localparam integer b145 = 5;
        for (m145 = 0; m145 < 16; m145 = m145 + 1) 
        begin: inbit145
            assign data_11[m145 + b145*16 + a5*28*16] = data_11_array[a5][b145][m145];
        end
    endgenerate
    generate 
        localparam integer b146 = 6;
        for (m146 = 0; m146 < 16; m146 = m146 + 1) 
        begin: inbit146
            assign data_11[m146 + b146*16 + a5*28*16] = data_11_array[a5][b146][m146];
        end
    endgenerate
    generate 
        localparam integer b147 = 7;
        for (m147 = 0; m147 < 16; m147 = m147 + 1) 
        begin: inbit147
            assign data_11[m147 + b147*16 + a5*28*16] = data_11_array[a5][b147][m147];
        end
    endgenerate
    generate 
        localparam integer b148 = 8;
        for (m148 = 0; m148 < 16; m148 = m148 + 1) 
        begin: inbit148
            assign data_11[m148 + b148*16 + a5*28*16] = data_11_array[a5][b148][m148];
        end
    endgenerate
    generate 
        localparam integer b149 = 9;
        for (m149 = 0; m149 < 16; m149 = m149 + 1) 
        begin: inbit149
            assign data_11[m149 + b149*16 + a5*28*16] = data_11_array[a5][b149][m149];
        end
    endgenerate
    generate 
        localparam integer b150 = 10;
        for (m150 = 0; m150 < 16; m150 = m150 + 1) 
        begin: inbit150
            assign data_11[m150 + b150*16 + a5*28*16] = data_11_array[a5][b150][m150];
        end
    endgenerate
    generate 
        localparam integer b151 = 11;
        for (m151 = 0; m151 < 16; m151 = m151 + 1) 
        begin: inbit151
            assign data_11[m151 + b151*16 + a5*28*16] = data_11_array[a5][b151][m151];
        end
    endgenerate
    generate 
        localparam integer b152 = 12;
        for (m152 = 0; m152 < 16; m152 = m152 + 1) 
        begin: inbit152
            assign data_11[m152 + b152*16 + a5*28*16] = data_11_array[a5][b152][m152];
        end
    endgenerate
    generate 
        localparam integer b153 = 13;
        for (m153 = 0; m153 < 16; m153 = m153 + 1) 
        begin: inbit153
            assign data_11[m153 + b153*16 + a5*28*16] = data_11_array[a5][b153][m153];
        end
    endgenerate
    generate 
        localparam integer b154 = 14;
        for (m154 = 0; m154 < 16; m154 = m154 + 1) 
        begin: inbit154
            assign data_11[m154 + b154*16 + a5*28*16] = data_11_array[a5][b154][m154];
        end
    endgenerate
    generate 
        localparam integer b155 = 15;
        for (m155 = 0; m155 < 16; m155 = m155 + 1) 
        begin: inbit155
            assign data_11[m155 + b155*16 + a5*28*16] = data_11_array[a5][b155][m155];
        end
    endgenerate
    generate 
        localparam integer b156 = 16;
        for (m156 = 0; m156 < 16; m156 = m156 + 1) 
        begin: inbit156
            assign data_11[m156 + b156*16 + a5*28*16] = data_11_array[a5][b156][m156];
        end
    endgenerate
    generate 
        localparam integer b157 = 17;
        for (m157 = 0; m157 < 16; m157 = m157 + 1) 
        begin: inbit157
            assign data_11[m157 + b157*16 + a5*28*16] = data_11_array[a5][b157][m157];
        end
    endgenerate
    generate 
        localparam integer b158 = 18;
        for (m158 = 0; m158 < 16; m158 = m158 + 1) 
        begin: inbit158
            assign data_11[m158 + b158*16 + a5*28*16] = data_11_array[a5][b158][m158];
        end
    endgenerate
    generate 
        localparam integer b159 = 19;
        for (m159 = 0; m159 < 16; m159 = m159 + 1) 
        begin: inbit159
            assign data_11[m159 + b159*16 + a5*28*16] = data_11_array[a5][b159][m159];
        end
    endgenerate
    generate 
        localparam integer b160 = 20;
        for (m160 = 0; m160 < 16; m160 = m160 + 1) 
        begin: inbit160
            assign data_11[m160 + b160*16 + a5*28*16] = data_11_array[a5][b160][m160];
        end
    endgenerate
    generate 
        localparam integer b161 = 21;
        for (m161 = 0; m161 < 16; m161 = m161 + 1) 
        begin: inbit161
            assign data_11[m161 + b161*16 + a5*28*16] = data_11_array[a5][b161][m161];
        end
    endgenerate
    generate 
        localparam integer b162 = 22;
        for (m162 = 0; m162 < 16; m162 = m162 + 1) 
        begin: inbit162
            assign data_11[m162 + b162*16 + a5*28*16] = data_11_array[a5][b162][m162];
        end
    endgenerate
    generate 
        localparam integer b163 = 23;
        for (m163 = 0; m163 < 16; m163 = m163 + 1) 
        begin: inbit163
            assign data_11[m163 + b163*16 + a5*28*16] = data_11_array[a5][b163][m163];
        end
    endgenerate
    generate 
        localparam integer b164 = 24;
        for (m164 = 0; m164 < 16; m164 = m164 + 1) 
        begin: inbit164
            assign data_11[m164 + b164*16 + a5*28*16] = data_11_array[a5][b164][m164];
        end
    endgenerate
    generate 
        localparam integer b165 = 25;
        for (m165 = 0; m165 < 16; m165 = m165 + 1) 
        begin: inbit165
            assign data_11[m165 + b165*16 + a5*28*16] = data_11_array[a5][b165][m165];
        end
    endgenerate
    generate 
        localparam integer b166 = 26;
        for (m166 = 0; m166 < 16; m166 = m166 + 1) 
        begin: inbit166
            assign data_11[m166 + b166*16 + a5*28*16] = data_11_array[a5][b166][m166];
        end
    endgenerate
    generate 
        localparam integer b167 = 27;
        for (m167 = 0; m167 < 16; m167 = m167 + 1) 
        begin: inbit167
            assign data_11[m167 + b167*16 + a5*28*16] = data_11_array[a5][b167][m167];
        end
    endgenerate
    localparam integer a6 = 6;
    generate 
        localparam integer b168 = 0;
        for (m168 = 0; m168 < 16; m168 = m168 + 1) 
        begin: inbit168
            assign data_11[m168 + b168*16 + a6*28*16] = data_11_array[a6][b168][m168];
        end
    endgenerate
    generate 
        localparam integer b169 = 1;
        for (m169 = 0; m169 < 16; m169 = m169 + 1) 
        begin: inbit169
            assign data_11[m169 + b169*16 + a6*28*16] = data_11_array[a6][b169][m169];
        end
    endgenerate
    generate 
        localparam integer b170 = 2;
        for (m170 = 0; m170 < 16; m170 = m170 + 1) 
        begin: inbit170
            assign data_11[m170 + b170*16 + a6*28*16] = data_11_array[a6][b170][m170];
        end
    endgenerate
    generate 
        localparam integer b171 = 3;
        for (m171 = 0; m171 < 16; m171 = m171 + 1) 
        begin: inbit171
            assign data_11[m171 + b171*16 + a6*28*16] = data_11_array[a6][b171][m171];
        end
    endgenerate
    generate 
        localparam integer b172 = 4;
        for (m172 = 0; m172 < 16; m172 = m172 + 1) 
        begin: inbit172
            assign data_11[m172 + b172*16 + a6*28*16] = data_11_array[a6][b172][m172];
        end
    endgenerate
    generate 
        localparam integer b173 = 5;
        for (m173 = 0; m173 < 16; m173 = m173 + 1) 
        begin: inbit173
            assign data_11[m173 + b173*16 + a6*28*16] = data_11_array[a6][b173][m173];
        end
    endgenerate
    generate 
        localparam integer b174 = 6;
        for (m174 = 0; m174 < 16; m174 = m174 + 1) 
        begin: inbit174
            assign data_11[m174 + b174*16 + a6*28*16] = data_11_array[a6][b174][m174];
        end
    endgenerate
    generate 
        localparam integer b175 = 7;
        for (m175 = 0; m175 < 16; m175 = m175 + 1) 
        begin: inbit175
            assign data_11[m175 + b175*16 + a6*28*16] = data_11_array[a6][b175][m175];
        end
    endgenerate
    generate 
        localparam integer b176 = 8;
        for (m176 = 0; m176 < 16; m176 = m176 + 1) 
        begin: inbit176
            assign data_11[m176 + b176*16 + a6*28*16] = data_11_array[a6][b176][m176];
        end
    endgenerate
    generate 
        localparam integer b177 = 9;
        for (m177 = 0; m177 < 16; m177 = m177 + 1) 
        begin: inbit177
            assign data_11[m177 + b177*16 + a6*28*16] = data_11_array[a6][b177][m177];
        end
    endgenerate
    generate 
        localparam integer b178 = 10;
        for (m178 = 0; m178 < 16; m178 = m178 + 1) 
        begin: inbit178
            assign data_11[m178 + b178*16 + a6*28*16] = data_11_array[a6][b178][m178];
        end
    endgenerate
    generate 
        localparam integer b179 = 11;
        for (m179 = 0; m179 < 16; m179 = m179 + 1) 
        begin: inbit179
            assign data_11[m179 + b179*16 + a6*28*16] = data_11_array[a6][b179][m179];
        end
    endgenerate
    generate 
        localparam integer b180 = 12;
        for (m180 = 0; m180 < 16; m180 = m180 + 1) 
        begin: inbit180
            assign data_11[m180 + b180*16 + a6*28*16] = data_11_array[a6][b180][m180];
        end
    endgenerate
    generate 
        localparam integer b181 = 13;
        for (m181 = 0; m181 < 16; m181 = m181 + 1) 
        begin: inbit181
            assign data_11[m181 + b181*16 + a6*28*16] = data_11_array[a6][b181][m181];
        end
    endgenerate
    generate 
        localparam integer b182 = 14;
        for (m182 = 0; m182 < 16; m182 = m182 + 1) 
        begin: inbit182
            assign data_11[m182 + b182*16 + a6*28*16] = data_11_array[a6][b182][m182];
        end
    endgenerate
    generate 
        localparam integer b183 = 15;
        for (m183 = 0; m183 < 16; m183 = m183 + 1) 
        begin: inbit183
            assign data_11[m183 + b183*16 + a6*28*16] = data_11_array[a6][b183][m183];
        end
    endgenerate
    generate 
        localparam integer b184 = 16;
        for (m184 = 0; m184 < 16; m184 = m184 + 1) 
        begin: inbit184
            assign data_11[m184 + b184*16 + a6*28*16] = data_11_array[a6][b184][m184];
        end
    endgenerate
    generate 
        localparam integer b185 = 17;
        for (m185 = 0; m185 < 16; m185 = m185 + 1) 
        begin: inbit185
            assign data_11[m185 + b185*16 + a6*28*16] = data_11_array[a6][b185][m185];
        end
    endgenerate
    generate 
        localparam integer b186 = 18;
        for (m186 = 0; m186 < 16; m186 = m186 + 1) 
        begin: inbit186
            assign data_11[m186 + b186*16 + a6*28*16] = data_11_array[a6][b186][m186];
        end
    endgenerate
    generate 
        localparam integer b187 = 19;
        for (m187 = 0; m187 < 16; m187 = m187 + 1) 
        begin: inbit187
            assign data_11[m187 + b187*16 + a6*28*16] = data_11_array[a6][b187][m187];
        end
    endgenerate
    generate 
        localparam integer b188 = 20;
        for (m188 = 0; m188 < 16; m188 = m188 + 1) 
        begin: inbit188
            assign data_11[m188 + b188*16 + a6*28*16] = data_11_array[a6][b188][m188];
        end
    endgenerate
    generate 
        localparam integer b189 = 21;
        for (m189 = 0; m189 < 16; m189 = m189 + 1) 
        begin: inbit189
            assign data_11[m189 + b189*16 + a6*28*16] = data_11_array[a6][b189][m189];
        end
    endgenerate
    generate 
        localparam integer b190 = 22;
        for (m190 = 0; m190 < 16; m190 = m190 + 1) 
        begin: inbit190
            assign data_11[m190 + b190*16 + a6*28*16] = data_11_array[a6][b190][m190];
        end
    endgenerate
    generate 
        localparam integer b191 = 23;
        for (m191 = 0; m191 < 16; m191 = m191 + 1) 
        begin: inbit191
            assign data_11[m191 + b191*16 + a6*28*16] = data_11_array[a6][b191][m191];
        end
    endgenerate
    generate 
        localparam integer b192 = 24;
        for (m192 = 0; m192 < 16; m192 = m192 + 1) 
        begin: inbit192
            assign data_11[m192 + b192*16 + a6*28*16] = data_11_array[a6][b192][m192];
        end
    endgenerate
    generate 
        localparam integer b193 = 25;
        for (m193 = 0; m193 < 16; m193 = m193 + 1) 
        begin: inbit193
            assign data_11[m193 + b193*16 + a6*28*16] = data_11_array[a6][b193][m193];
        end
    endgenerate
    generate 
        localparam integer b194 = 26;
        for (m194 = 0; m194 < 16; m194 = m194 + 1) 
        begin: inbit194
            assign data_11[m194 + b194*16 + a6*28*16] = data_11_array[a6][b194][m194];
        end
    endgenerate
    generate 
        localparam integer b195 = 27;
        for (m195 = 0; m195 < 16; m195 = m195 + 1) 
        begin: inbit195
            assign data_11[m195 + b195*16 + a6*28*16] = data_11_array[a6][b195][m195];
        end
    endgenerate
    localparam integer a7 = 7;
    generate 
        localparam integer b196 = 0;
        for (m196 = 0; m196 < 16; m196 = m196 + 1) 
        begin: inbit196
            assign data_11[m196 + b196*16 + a7*28*16] = data_11_array[a7][b196][m196];
        end
    endgenerate
    generate 
        localparam integer b197 = 1;
        for (m197 = 0; m197 < 16; m197 = m197 + 1) 
        begin: inbit197
            assign data_11[m197 + b197*16 + a7*28*16] = data_11_array[a7][b197][m197];
        end
    endgenerate
    generate 
        localparam integer b198 = 2;
        for (m198 = 0; m198 < 16; m198 = m198 + 1) 
        begin: inbit198
            assign data_11[m198 + b198*16 + a7*28*16] = data_11_array[a7][b198][m198];
        end
    endgenerate
    generate 
        localparam integer b199 = 3;
        for (m199 = 0; m199 < 16; m199 = m199 + 1) 
        begin: inbit199
            assign data_11[m199 + b199*16 + a7*28*16] = data_11_array[a7][b199][m199];
        end
    endgenerate
    generate 
        localparam integer b200 = 4;
        for (m200 = 0; m200 < 16; m200 = m200 + 1) 
        begin: inbit200
            assign data_11[m200 + b200*16 + a7*28*16] = data_11_array[a7][b200][m200];
        end
    endgenerate
    generate 
        localparam integer b201 = 5;
        for (m201 = 0; m201 < 16; m201 = m201 + 1) 
        begin: inbit201
            assign data_11[m201 + b201*16 + a7*28*16] = data_11_array[a7][b201][m201];
        end
    endgenerate
    generate 
        localparam integer b202 = 6;
        for (m202 = 0; m202 < 16; m202 = m202 + 1) 
        begin: inbit202
            assign data_11[m202 + b202*16 + a7*28*16] = data_11_array[a7][b202][m202];
        end
    endgenerate
    generate 
        localparam integer b203 = 7;
        for (m203 = 0; m203 < 16; m203 = m203 + 1) 
        begin: inbit203
            assign data_11[m203 + b203*16 + a7*28*16] = data_11_array[a7][b203][m203];
        end
    endgenerate
    generate 
        localparam integer b204 = 8;
        for (m204 = 0; m204 < 16; m204 = m204 + 1) 
        begin: inbit204
            assign data_11[m204 + b204*16 + a7*28*16] = data_11_array[a7][b204][m204];
        end
    endgenerate
    generate 
        localparam integer b205 = 9;
        for (m205 = 0; m205 < 16; m205 = m205 + 1) 
        begin: inbit205
            assign data_11[m205 + b205*16 + a7*28*16] = data_11_array[a7][b205][m205];
        end
    endgenerate
    generate 
        localparam integer b206 = 10;
        for (m206 = 0; m206 < 16; m206 = m206 + 1) 
        begin: inbit206
            assign data_11[m206 + b206*16 + a7*28*16] = data_11_array[a7][b206][m206];
        end
    endgenerate
    generate 
        localparam integer b207 = 11;
        for (m207 = 0; m207 < 16; m207 = m207 + 1) 
        begin: inbit207
            assign data_11[m207 + b207*16 + a7*28*16] = data_11_array[a7][b207][m207];
        end
    endgenerate
    generate 
        localparam integer b208 = 12;
        for (m208 = 0; m208 < 16; m208 = m208 + 1) 
        begin: inbit208
            assign data_11[m208 + b208*16 + a7*28*16] = data_11_array[a7][b208][m208];
        end
    endgenerate
    generate 
        localparam integer b209 = 13;
        for (m209 = 0; m209 < 16; m209 = m209 + 1) 
        begin: inbit209
            assign data_11[m209 + b209*16 + a7*28*16] = data_11_array[a7][b209][m209];
        end
    endgenerate
    generate 
        localparam integer b210 = 14;
        for (m210 = 0; m210 < 16; m210 = m210 + 1) 
        begin: inbit210
            assign data_11[m210 + b210*16 + a7*28*16] = data_11_array[a7][b210][m210];
        end
    endgenerate
    generate 
        localparam integer b211 = 15;
        for (m211 = 0; m211 < 16; m211 = m211 + 1) 
        begin: inbit211
            assign data_11[m211 + b211*16 + a7*28*16] = data_11_array[a7][b211][m211];
        end
    endgenerate
    generate 
        localparam integer b212 = 16;
        for (m212 = 0; m212 < 16; m212 = m212 + 1) 
        begin: inbit212
            assign data_11[m212 + b212*16 + a7*28*16] = data_11_array[a7][b212][m212];
        end
    endgenerate
    generate 
        localparam integer b213 = 17;
        for (m213 = 0; m213 < 16; m213 = m213 + 1) 
        begin: inbit213
            assign data_11[m213 + b213*16 + a7*28*16] = data_11_array[a7][b213][m213];
        end
    endgenerate
    generate 
        localparam integer b214 = 18;
        for (m214 = 0; m214 < 16; m214 = m214 + 1) 
        begin: inbit214
            assign data_11[m214 + b214*16 + a7*28*16] = data_11_array[a7][b214][m214];
        end
    endgenerate
    generate 
        localparam integer b215 = 19;
        for (m215 = 0; m215 < 16; m215 = m215 + 1) 
        begin: inbit215
            assign data_11[m215 + b215*16 + a7*28*16] = data_11_array[a7][b215][m215];
        end
    endgenerate
    generate 
        localparam integer b216 = 20;
        for (m216 = 0; m216 < 16; m216 = m216 + 1) 
        begin: inbit216
            assign data_11[m216 + b216*16 + a7*28*16] = data_11_array[a7][b216][m216];
        end
    endgenerate
    generate 
        localparam integer b217 = 21;
        for (m217 = 0; m217 < 16; m217 = m217 + 1) 
        begin: inbit217
            assign data_11[m217 + b217*16 + a7*28*16] = data_11_array[a7][b217][m217];
        end
    endgenerate
    generate 
        localparam integer b218 = 22;
        for (m218 = 0; m218 < 16; m218 = m218 + 1) 
        begin: inbit218
            assign data_11[m218 + b218*16 + a7*28*16] = data_11_array[a7][b218][m218];
        end
    endgenerate
    generate 
        localparam integer b219 = 23;
        for (m219 = 0; m219 < 16; m219 = m219 + 1) 
        begin: inbit219
            assign data_11[m219 + b219*16 + a7*28*16] = data_11_array[a7][b219][m219];
        end
    endgenerate
    generate 
        localparam integer b220 = 24;
        for (m220 = 0; m220 < 16; m220 = m220 + 1) 
        begin: inbit220
            assign data_11[m220 + b220*16 + a7*28*16] = data_11_array[a7][b220][m220];
        end
    endgenerate
    generate 
        localparam integer b221 = 25;
        for (m221 = 0; m221 < 16; m221 = m221 + 1) 
        begin: inbit221
            assign data_11[m221 + b221*16 + a7*28*16] = data_11_array[a7][b221][m221];
        end
    endgenerate
    generate 
        localparam integer b222 = 26;
        for (m222 = 0; m222 < 16; m222 = m222 + 1) 
        begin: inbit222
            assign data_11[m222 + b222*16 + a7*28*16] = data_11_array[a7][b222][m222];
        end
    endgenerate
    generate 
        localparam integer b223 = 27;
        for (m223 = 0; m223 < 16; m223 = m223 + 1) 
        begin: inbit223
            assign data_11[m223 + b223*16 + a7*28*16] = data_11_array[a7][b223][m223];
        end
    endgenerate
    localparam integer a8 = 8;
    generate 
        localparam integer b224 = 0;
        for (m224 = 0; m224 < 16; m224 = m224 + 1) 
        begin: inbit224
            assign data_11[m224 + b224*16 + a8*28*16] = data_11_array[a8][b224][m224];
        end
    endgenerate
    generate 
        localparam integer b225 = 1;
        for (m225 = 0; m225 < 16; m225 = m225 + 1) 
        begin: inbit225
            assign data_11[m225 + b225*16 + a8*28*16] = data_11_array[a8][b225][m225];
        end
    endgenerate
    generate 
        localparam integer b226 = 2;
        for (m226 = 0; m226 < 16; m226 = m226 + 1) 
        begin: inbit226
            assign data_11[m226 + b226*16 + a8*28*16] = data_11_array[a8][b226][m226];
        end
    endgenerate
    generate 
        localparam integer b227 = 3;
        for (m227 = 0; m227 < 16; m227 = m227 + 1) 
        begin: inbit227
            assign data_11[m227 + b227*16 + a8*28*16] = data_11_array[a8][b227][m227];
        end
    endgenerate
    generate 
        localparam integer b228 = 4;
        for (m228 = 0; m228 < 16; m228 = m228 + 1) 
        begin: inbit228
            assign data_11[m228 + b228*16 + a8*28*16] = data_11_array[a8][b228][m228];
        end
    endgenerate
    generate 
        localparam integer b229 = 5;
        for (m229 = 0; m229 < 16; m229 = m229 + 1) 
        begin: inbit229
            assign data_11[m229 + b229*16 + a8*28*16] = data_11_array[a8][b229][m229];
        end
    endgenerate
    generate 
        localparam integer b230 = 6;
        for (m230 = 0; m230 < 16; m230 = m230 + 1) 
        begin: inbit230
            assign data_11[m230 + b230*16 + a8*28*16] = data_11_array[a8][b230][m230];
        end
    endgenerate
    generate 
        localparam integer b231 = 7;
        for (m231 = 0; m231 < 16; m231 = m231 + 1) 
        begin: inbit231
            assign data_11[m231 + b231*16 + a8*28*16] = data_11_array[a8][b231][m231];
        end
    endgenerate
    generate 
        localparam integer b232 = 8;
        for (m232 = 0; m232 < 16; m232 = m232 + 1) 
        begin: inbit232
            assign data_11[m232 + b232*16 + a8*28*16] = data_11_array[a8][b232][m232];
        end
    endgenerate
    generate 
        localparam integer b233 = 9;
        for (m233 = 0; m233 < 16; m233 = m233 + 1) 
        begin: inbit233
            assign data_11[m233 + b233*16 + a8*28*16] = data_11_array[a8][b233][m233];
        end
    endgenerate
    generate 
        localparam integer b234 = 10;
        for (m234 = 0; m234 < 16; m234 = m234 + 1) 
        begin: inbit234
            assign data_11[m234 + b234*16 + a8*28*16] = data_11_array[a8][b234][m234];
        end
    endgenerate
    generate 
        localparam integer b235 = 11;
        for (m235 = 0; m235 < 16; m235 = m235 + 1) 
        begin: inbit235
            assign data_11[m235 + b235*16 + a8*28*16] = data_11_array[a8][b235][m235];
        end
    endgenerate
    generate 
        localparam integer b236 = 12;
        for (m236 = 0; m236 < 16; m236 = m236 + 1) 
        begin: inbit236
            assign data_11[m236 + b236*16 + a8*28*16] = data_11_array[a8][b236][m236];
        end
    endgenerate
    generate 
        localparam integer b237 = 13;
        for (m237 = 0; m237 < 16; m237 = m237 + 1) 
        begin: inbit237
            assign data_11[m237 + b237*16 + a8*28*16] = data_11_array[a8][b237][m237];
        end
    endgenerate
    generate 
        localparam integer b238 = 14;
        for (m238 = 0; m238 < 16; m238 = m238 + 1) 
        begin: inbit238
            assign data_11[m238 + b238*16 + a8*28*16] = data_11_array[a8][b238][m238];
        end
    endgenerate
    generate 
        localparam integer b239 = 15;
        for (m239 = 0; m239 < 16; m239 = m239 + 1) 
        begin: inbit239
            assign data_11[m239 + b239*16 + a8*28*16] = data_11_array[a8][b239][m239];
        end
    endgenerate
    generate 
        localparam integer b240 = 16;
        for (m240 = 0; m240 < 16; m240 = m240 + 1) 
        begin: inbit240
            assign data_11[m240 + b240*16 + a8*28*16] = data_11_array[a8][b240][m240];
        end
    endgenerate
    generate 
        localparam integer b241 = 17;
        for (m241 = 0; m241 < 16; m241 = m241 + 1) 
        begin: inbit241
            assign data_11[m241 + b241*16 + a8*28*16] = data_11_array[a8][b241][m241];
        end
    endgenerate
    generate 
        localparam integer b242 = 18;
        for (m242 = 0; m242 < 16; m242 = m242 + 1) 
        begin: inbit242
            assign data_11[m242 + b242*16 + a8*28*16] = data_11_array[a8][b242][m242];
        end
    endgenerate
    generate 
        localparam integer b243 = 19;
        for (m243 = 0; m243 < 16; m243 = m243 + 1) 
        begin: inbit243
            assign data_11[m243 + b243*16 + a8*28*16] = data_11_array[a8][b243][m243];
        end
    endgenerate
    generate 
        localparam integer b244 = 20;
        for (m244 = 0; m244 < 16; m244 = m244 + 1) 
        begin: inbit244
            assign data_11[m244 + b244*16 + a8*28*16] = data_11_array[a8][b244][m244];
        end
    endgenerate
    generate 
        localparam integer b245 = 21;
        for (m245 = 0; m245 < 16; m245 = m245 + 1) 
        begin: inbit245
            assign data_11[m245 + b245*16 + a8*28*16] = data_11_array[a8][b245][m245];
        end
    endgenerate
    generate 
        localparam integer b246 = 22;
        for (m246 = 0; m246 < 16; m246 = m246 + 1) 
        begin: inbit246
            assign data_11[m246 + b246*16 + a8*28*16] = data_11_array[a8][b246][m246];
        end
    endgenerate
    generate 
        localparam integer b247 = 23;
        for (m247 = 0; m247 < 16; m247 = m247 + 1) 
        begin: inbit247
            assign data_11[m247 + b247*16 + a8*28*16] = data_11_array[a8][b247][m247];
        end
    endgenerate
    generate 
        localparam integer b248 = 24;
        for (m248 = 0; m248 < 16; m248 = m248 + 1) 
        begin: inbit248
            assign data_11[m248 + b248*16 + a8*28*16] = data_11_array[a8][b248][m248];
        end
    endgenerate
    generate 
        localparam integer b249 = 25;
        for (m249 = 0; m249 < 16; m249 = m249 + 1) 
        begin: inbit249
            assign data_11[m249 + b249*16 + a8*28*16] = data_11_array[a8][b249][m249];
        end
    endgenerate
    generate 
        localparam integer b250 = 26;
        for (m250 = 0; m250 < 16; m250 = m250 + 1) 
        begin: inbit250
            assign data_11[m250 + b250*16 + a8*28*16] = data_11_array[a8][b250][m250];
        end
    endgenerate
    generate 
        localparam integer b251 = 27;
        for (m251 = 0; m251 < 16; m251 = m251 + 1) 
        begin: inbit251
            assign data_11[m251 + b251*16 + a8*28*16] = data_11_array[a8][b251][m251];
        end
    endgenerate
    localparam integer a9 = 9;
    generate 
        localparam integer b252 = 0;
        for (m252 = 0; m252 < 16; m252 = m252 + 1) 
        begin: inbit252
            assign data_11[m252 + b252*16 + a9*28*16] = data_11_array[a9][b252][m252];
        end
    endgenerate
    generate 
        localparam integer b253 = 1;
        for (m253 = 0; m253 < 16; m253 = m253 + 1) 
        begin: inbit253
            assign data_11[m253 + b253*16 + a9*28*16] = data_11_array[a9][b253][m253];
        end
    endgenerate
    generate 
        localparam integer b254 = 2;
        for (m254 = 0; m254 < 16; m254 = m254 + 1) 
        begin: inbit254
            assign data_11[m254 + b254*16 + a9*28*16] = data_11_array[a9][b254][m254];
        end
    endgenerate
    generate 
        localparam integer b255 = 3;
        for (m255 = 0; m255 < 16; m255 = m255 + 1) 
        begin: inbit255
            assign data_11[m255 + b255*16 + a9*28*16] = data_11_array[a9][b255][m255];
        end
    endgenerate
    generate 
        localparam integer b256 = 4;
        for (m256 = 0; m256 < 16; m256 = m256 + 1) 
        begin: inbit256
            assign data_11[m256 + b256*16 + a9*28*16] = data_11_array[a9][b256][m256];
        end
    endgenerate
    generate 
        localparam integer b257 = 5;
        for (m257 = 0; m257 < 16; m257 = m257 + 1) 
        begin: inbit257
            assign data_11[m257 + b257*16 + a9*28*16] = data_11_array[a9][b257][m257];
        end
    endgenerate
    generate 
        localparam integer b258 = 6;
        for (m258 = 0; m258 < 16; m258 = m258 + 1) 
        begin: inbit258
            assign data_11[m258 + b258*16 + a9*28*16] = data_11_array[a9][b258][m258];
        end
    endgenerate
    generate 
        localparam integer b259 = 7;
        for (m259 = 0; m259 < 16; m259 = m259 + 1) 
        begin: inbit259
            assign data_11[m259 + b259*16 + a9*28*16] = data_11_array[a9][b259][m259];
        end
    endgenerate
    generate 
        localparam integer b260 = 8;
        for (m260 = 0; m260 < 16; m260 = m260 + 1) 
        begin: inbit260
            assign data_11[m260 + b260*16 + a9*28*16] = data_11_array[a9][b260][m260];
        end
    endgenerate
    generate 
        localparam integer b261 = 9;
        for (m261 = 0; m261 < 16; m261 = m261 + 1) 
        begin: inbit261
            assign data_11[m261 + b261*16 + a9*28*16] = data_11_array[a9][b261][m261];
        end
    endgenerate
    generate 
        localparam integer b262 = 10;
        for (m262 = 0; m262 < 16; m262 = m262 + 1) 
        begin: inbit262
            assign data_11[m262 + b262*16 + a9*28*16] = data_11_array[a9][b262][m262];
        end
    endgenerate
    generate 
        localparam integer b263 = 11;
        for (m263 = 0; m263 < 16; m263 = m263 + 1) 
        begin: inbit263
            assign data_11[m263 + b263*16 + a9*28*16] = data_11_array[a9][b263][m263];
        end
    endgenerate
    generate 
        localparam integer b264 = 12;
        for (m264 = 0; m264 < 16; m264 = m264 + 1) 
        begin: inbit264
            assign data_11[m264 + b264*16 + a9*28*16] = data_11_array[a9][b264][m264];
        end
    endgenerate
    generate 
        localparam integer b265 = 13;
        for (m265 = 0; m265 < 16; m265 = m265 + 1) 
        begin: inbit265
            assign data_11[m265 + b265*16 + a9*28*16] = data_11_array[a9][b265][m265];
        end
    endgenerate
    generate 
        localparam integer b266 = 14;
        for (m266 = 0; m266 < 16; m266 = m266 + 1) 
        begin: inbit266
            assign data_11[m266 + b266*16 + a9*28*16] = data_11_array[a9][b266][m266];
        end
    endgenerate
    generate 
        localparam integer b267 = 15;
        for (m267 = 0; m267 < 16; m267 = m267 + 1) 
        begin: inbit267
            assign data_11[m267 + b267*16 + a9*28*16] = data_11_array[a9][b267][m267];
        end
    endgenerate
    generate 
        localparam integer b268 = 16;
        for (m268 = 0; m268 < 16; m268 = m268 + 1) 
        begin: inbit268
            assign data_11[m268 + b268*16 + a9*28*16] = data_11_array[a9][b268][m268];
        end
    endgenerate
    generate 
        localparam integer b269 = 17;
        for (m269 = 0; m269 < 16; m269 = m269 + 1) 
        begin: inbit269
            assign data_11[m269 + b269*16 + a9*28*16] = data_11_array[a9][b269][m269];
        end
    endgenerate
    generate 
        localparam integer b270 = 18;
        for (m270 = 0; m270 < 16; m270 = m270 + 1) 
        begin: inbit270
            assign data_11[m270 + b270*16 + a9*28*16] = data_11_array[a9][b270][m270];
        end
    endgenerate
    generate 
        localparam integer b271 = 19;
        for (m271 = 0; m271 < 16; m271 = m271 + 1) 
        begin: inbit271
            assign data_11[m271 + b271*16 + a9*28*16] = data_11_array[a9][b271][m271];
        end
    endgenerate
    generate 
        localparam integer b272 = 20;
        for (m272 = 0; m272 < 16; m272 = m272 + 1) 
        begin: inbit272
            assign data_11[m272 + b272*16 + a9*28*16] = data_11_array[a9][b272][m272];
        end
    endgenerate
    generate 
        localparam integer b273 = 21;
        for (m273 = 0; m273 < 16; m273 = m273 + 1) 
        begin: inbit273
            assign data_11[m273 + b273*16 + a9*28*16] = data_11_array[a9][b273][m273];
        end
    endgenerate
    generate 
        localparam integer b274 = 22;
        for (m274 = 0; m274 < 16; m274 = m274 + 1) 
        begin: inbit274
            assign data_11[m274 + b274*16 + a9*28*16] = data_11_array[a9][b274][m274];
        end
    endgenerate
    generate 
        localparam integer b275 = 23;
        for (m275 = 0; m275 < 16; m275 = m275 + 1) 
        begin: inbit275
            assign data_11[m275 + b275*16 + a9*28*16] = data_11_array[a9][b275][m275];
        end
    endgenerate
    generate 
        localparam integer b276 = 24;
        for (m276 = 0; m276 < 16; m276 = m276 + 1) 
        begin: inbit276
            assign data_11[m276 + b276*16 + a9*28*16] = data_11_array[a9][b276][m276];
        end
    endgenerate
    generate 
        localparam integer b277 = 25;
        for (m277 = 0; m277 < 16; m277 = m277 + 1) 
        begin: inbit277
            assign data_11[m277 + b277*16 + a9*28*16] = data_11_array[a9][b277][m277];
        end
    endgenerate
    generate 
        localparam integer b278 = 26;
        for (m278 = 0; m278 < 16; m278 = m278 + 1) 
        begin: inbit278
            assign data_11[m278 + b278*16 + a9*28*16] = data_11_array[a9][b278][m278];
        end
    endgenerate
    generate 
        localparam integer b279 = 27;
        for (m279 = 0; m279 < 16; m279 = m279 + 1) 
        begin: inbit279
            assign data_11[m279 + b279*16 + a9*28*16] = data_11_array[a9][b279][m279];
        end
    endgenerate
    localparam integer a10 = 10;
    generate 
        localparam integer b280 = 0;
        for (m280 = 0; m280 < 16; m280 = m280 + 1) 
        begin: inbit280
            assign data_11[m280 + b280*16 + a10*28*16] = data_11_array[a10][b280][m280];
        end
    endgenerate
    generate 
        localparam integer b281 = 1;
        for (m281 = 0; m281 < 16; m281 = m281 + 1) 
        begin: inbit281
            assign data_11[m281 + b281*16 + a10*28*16] = data_11_array[a10][b281][m281];
        end
    endgenerate
    generate 
        localparam integer b282 = 2;
        for (m282 = 0; m282 < 16; m282 = m282 + 1) 
        begin: inbit282
            assign data_11[m282 + b282*16 + a10*28*16] = data_11_array[a10][b282][m282];
        end
    endgenerate
    generate 
        localparam integer b283 = 3;
        for (m283 = 0; m283 < 16; m283 = m283 + 1) 
        begin: inbit283
            assign data_11[m283 + b283*16 + a10*28*16] = data_11_array[a10][b283][m283];
        end
    endgenerate
    generate 
        localparam integer b284 = 4;
        for (m284 = 0; m284 < 16; m284 = m284 + 1) 
        begin: inbit284
            assign data_11[m284 + b284*16 + a10*28*16] = data_11_array[a10][b284][m284];
        end
    endgenerate
    generate 
        localparam integer b285 = 5;
        for (m285 = 0; m285 < 16; m285 = m285 + 1) 
        begin: inbit285
            assign data_11[m285 + b285*16 + a10*28*16] = data_11_array[a10][b285][m285];
        end
    endgenerate
    generate 
        localparam integer b286 = 6;
        for (m286 = 0; m286 < 16; m286 = m286 + 1) 
        begin: inbit286
            assign data_11[m286 + b286*16 + a10*28*16] = data_11_array[a10][b286][m286];
        end
    endgenerate
    generate 
        localparam integer b287 = 7;
        for (m287 = 0; m287 < 16; m287 = m287 + 1) 
        begin: inbit287
            assign data_11[m287 + b287*16 + a10*28*16] = data_11_array[a10][b287][m287];
        end
    endgenerate
    generate 
        localparam integer b288 = 8;
        for (m288 = 0; m288 < 16; m288 = m288 + 1) 
        begin: inbit288
            assign data_11[m288 + b288*16 + a10*28*16] = data_11_array[a10][b288][m288];
        end
    endgenerate
    generate 
        localparam integer b289 = 9;
        for (m289 = 0; m289 < 16; m289 = m289 + 1) 
        begin: inbit289
            assign data_11[m289 + b289*16 + a10*28*16] = data_11_array[a10][b289][m289];
        end
    endgenerate
    generate 
        localparam integer b290 = 10;
        for (m290 = 0; m290 < 16; m290 = m290 + 1) 
        begin: inbit290
            assign data_11[m290 + b290*16 + a10*28*16] = data_11_array[a10][b290][m290];
        end
    endgenerate
    generate 
        localparam integer b291 = 11;
        for (m291 = 0; m291 < 16; m291 = m291 + 1) 
        begin: inbit291
            assign data_11[m291 + b291*16 + a10*28*16] = data_11_array[a10][b291][m291];
        end
    endgenerate
    generate 
        localparam integer b292 = 12;
        for (m292 = 0; m292 < 16; m292 = m292 + 1) 
        begin: inbit292
            assign data_11[m292 + b292*16 + a10*28*16] = data_11_array[a10][b292][m292];
        end
    endgenerate
    generate 
        localparam integer b293 = 13;
        for (m293 = 0; m293 < 16; m293 = m293 + 1) 
        begin: inbit293
            assign data_11[m293 + b293*16 + a10*28*16] = data_11_array[a10][b293][m293];
        end
    endgenerate
    generate 
        localparam integer b294 = 14;
        for (m294 = 0; m294 < 16; m294 = m294 + 1) 
        begin: inbit294
            assign data_11[m294 + b294*16 + a10*28*16] = data_11_array[a10][b294][m294];
        end
    endgenerate
    generate 
        localparam integer b295 = 15;
        for (m295 = 0; m295 < 16; m295 = m295 + 1) 
        begin: inbit295
            assign data_11[m295 + b295*16 + a10*28*16] = data_11_array[a10][b295][m295];
        end
    endgenerate
    generate 
        localparam integer b296 = 16;
        for (m296 = 0; m296 < 16; m296 = m296 + 1) 
        begin: inbit296
            assign data_11[m296 + b296*16 + a10*28*16] = data_11_array[a10][b296][m296];
        end
    endgenerate
    generate 
        localparam integer b297 = 17;
        for (m297 = 0; m297 < 16; m297 = m297 + 1) 
        begin: inbit297
            assign data_11[m297 + b297*16 + a10*28*16] = data_11_array[a10][b297][m297];
        end
    endgenerate
    generate 
        localparam integer b298 = 18;
        for (m298 = 0; m298 < 16; m298 = m298 + 1) 
        begin: inbit298
            assign data_11[m298 + b298*16 + a10*28*16] = data_11_array[a10][b298][m298];
        end
    endgenerate
    generate 
        localparam integer b299 = 19;
        for (m299 = 0; m299 < 16; m299 = m299 + 1) 
        begin: inbit299
            assign data_11[m299 + b299*16 + a10*28*16] = data_11_array[a10][b299][m299];
        end
    endgenerate
    generate 
        localparam integer b300 = 20;
        for (m300 = 0; m300 < 16; m300 = m300 + 1) 
        begin: inbit300
            assign data_11[m300 + b300*16 + a10*28*16] = data_11_array[a10][b300][m300];
        end
    endgenerate
    generate 
        localparam integer b301 = 21;
        for (m301 = 0; m301 < 16; m301 = m301 + 1) 
        begin: inbit301
            assign data_11[m301 + b301*16 + a10*28*16] = data_11_array[a10][b301][m301];
        end
    endgenerate
    generate 
        localparam integer b302 = 22;
        for (m302 = 0; m302 < 16; m302 = m302 + 1) 
        begin: inbit302
            assign data_11[m302 + b302*16 + a10*28*16] = data_11_array[a10][b302][m302];
        end
    endgenerate
    generate 
        localparam integer b303 = 23;
        for (m303 = 0; m303 < 16; m303 = m303 + 1) 
        begin: inbit303
            assign data_11[m303 + b303*16 + a10*28*16] = data_11_array[a10][b303][m303];
        end
    endgenerate
    generate 
        localparam integer b304 = 24;
        for (m304 = 0; m304 < 16; m304 = m304 + 1) 
        begin: inbit304
            assign data_11[m304 + b304*16 + a10*28*16] = data_11_array[a10][b304][m304];
        end
    endgenerate
    generate 
        localparam integer b305 = 25;
        for (m305 = 0; m305 < 16; m305 = m305 + 1) 
        begin: inbit305
            assign data_11[m305 + b305*16 + a10*28*16] = data_11_array[a10][b305][m305];
        end
    endgenerate
    generate 
        localparam integer b306 = 26;
        for (m306 = 0; m306 < 16; m306 = m306 + 1) 
        begin: inbit306
            assign data_11[m306 + b306*16 + a10*28*16] = data_11_array[a10][b306][m306];
        end
    endgenerate
    generate 
        localparam integer b307 = 27;
        for (m307 = 0; m307 < 16; m307 = m307 + 1) 
        begin: inbit307
            assign data_11[m307 + b307*16 + a10*28*16] = data_11_array[a10][b307][m307];
        end
    endgenerate
    localparam integer a11 = 11;
    generate 
        localparam integer b308 = 0;
        for (m308 = 0; m308 < 16; m308 = m308 + 1) 
        begin: inbit308
            assign data_11[m308 + b308*16 + a11*28*16] = data_11_array[a11][b308][m308];
        end
    endgenerate
    generate 
        localparam integer b309 = 1;
        for (m309 = 0; m309 < 16; m309 = m309 + 1) 
        begin: inbit309
            assign data_11[m309 + b309*16 + a11*28*16] = data_11_array[a11][b309][m309];
        end
    endgenerate
    generate 
        localparam integer b310 = 2;
        for (m310 = 0; m310 < 16; m310 = m310 + 1) 
        begin: inbit310
            assign data_11[m310 + b310*16 + a11*28*16] = data_11_array[a11][b310][m310];
        end
    endgenerate
    generate 
        localparam integer b311 = 3;
        for (m311 = 0; m311 < 16; m311 = m311 + 1) 
        begin: inbit311
            assign data_11[m311 + b311*16 + a11*28*16] = data_11_array[a11][b311][m311];
        end
    endgenerate
    generate 
        localparam integer b312 = 4;
        for (m312 = 0; m312 < 16; m312 = m312 + 1) 
        begin: inbit312
            assign data_11[m312 + b312*16 + a11*28*16] = data_11_array[a11][b312][m312];
        end
    endgenerate
    generate 
        localparam integer b313 = 5;
        for (m313 = 0; m313 < 16; m313 = m313 + 1) 
        begin: inbit313
            assign data_11[m313 + b313*16 + a11*28*16] = data_11_array[a11][b313][m313];
        end
    endgenerate
    generate 
        localparam integer b314 = 6;
        for (m314 = 0; m314 < 16; m314 = m314 + 1) 
        begin: inbit314
            assign data_11[m314 + b314*16 + a11*28*16] = data_11_array[a11][b314][m314];
        end
    endgenerate
    generate 
        localparam integer b315 = 7;
        for (m315 = 0; m315 < 16; m315 = m315 + 1) 
        begin: inbit315
            assign data_11[m315 + b315*16 + a11*28*16] = data_11_array[a11][b315][m315];
        end
    endgenerate
    generate 
        localparam integer b316 = 8;
        for (m316 = 0; m316 < 16; m316 = m316 + 1) 
        begin: inbit316
            assign data_11[m316 + b316*16 + a11*28*16] = data_11_array[a11][b316][m316];
        end
    endgenerate
    generate 
        localparam integer b317 = 9;
        for (m317 = 0; m317 < 16; m317 = m317 + 1) 
        begin: inbit317
            assign data_11[m317 + b317*16 + a11*28*16] = data_11_array[a11][b317][m317];
        end
    endgenerate
    generate 
        localparam integer b318 = 10;
        for (m318 = 0; m318 < 16; m318 = m318 + 1) 
        begin: inbit318
            assign data_11[m318 + b318*16 + a11*28*16] = data_11_array[a11][b318][m318];
        end
    endgenerate
    generate 
        localparam integer b319 = 11;
        for (m319 = 0; m319 < 16; m319 = m319 + 1) 
        begin: inbit319
            assign data_11[m319 + b319*16 + a11*28*16] = data_11_array[a11][b319][m319];
        end
    endgenerate
    generate 
        localparam integer b320 = 12;
        for (m320 = 0; m320 < 16; m320 = m320 + 1) 
        begin: inbit320
            assign data_11[m320 + b320*16 + a11*28*16] = data_11_array[a11][b320][m320];
        end
    endgenerate
    generate 
        localparam integer b321 = 13;
        for (m321 = 0; m321 < 16; m321 = m321 + 1) 
        begin: inbit321
            assign data_11[m321 + b321*16 + a11*28*16] = data_11_array[a11][b321][m321];
        end
    endgenerate
    generate 
        localparam integer b322 = 14;
        for (m322 = 0; m322 < 16; m322 = m322 + 1) 
        begin: inbit322
            assign data_11[m322 + b322*16 + a11*28*16] = data_11_array[a11][b322][m322];
        end
    endgenerate
    generate 
        localparam integer b323 = 15;
        for (m323 = 0; m323 < 16; m323 = m323 + 1) 
        begin: inbit323
            assign data_11[m323 + b323*16 + a11*28*16] = data_11_array[a11][b323][m323];
        end
    endgenerate
    generate 
        localparam integer b324 = 16;
        for (m324 = 0; m324 < 16; m324 = m324 + 1) 
        begin: inbit324
            assign data_11[m324 + b324*16 + a11*28*16] = data_11_array[a11][b324][m324];
        end
    endgenerate
    generate 
        localparam integer b325 = 17;
        for (m325 = 0; m325 < 16; m325 = m325 + 1) 
        begin: inbit325
            assign data_11[m325 + b325*16 + a11*28*16] = data_11_array[a11][b325][m325];
        end
    endgenerate
    generate 
        localparam integer b326 = 18;
        for (m326 = 0; m326 < 16; m326 = m326 + 1) 
        begin: inbit326
            assign data_11[m326 + b326*16 + a11*28*16] = data_11_array[a11][b326][m326];
        end
    endgenerate
    generate 
        localparam integer b327 = 19;
        for (m327 = 0; m327 < 16; m327 = m327 + 1) 
        begin: inbit327
            assign data_11[m327 + b327*16 + a11*28*16] = data_11_array[a11][b327][m327];
        end
    endgenerate
    generate 
        localparam integer b328 = 20;
        for (m328 = 0; m328 < 16; m328 = m328 + 1) 
        begin: inbit328
            assign data_11[m328 + b328*16 + a11*28*16] = data_11_array[a11][b328][m328];
        end
    endgenerate
    generate 
        localparam integer b329 = 21;
        for (m329 = 0; m329 < 16; m329 = m329 + 1) 
        begin: inbit329
            assign data_11[m329 + b329*16 + a11*28*16] = data_11_array[a11][b329][m329];
        end
    endgenerate
    generate 
        localparam integer b330 = 22;
        for (m330 = 0; m330 < 16; m330 = m330 + 1) 
        begin: inbit330
            assign data_11[m330 + b330*16 + a11*28*16] = data_11_array[a11][b330][m330];
        end
    endgenerate
    generate 
        localparam integer b331 = 23;
        for (m331 = 0; m331 < 16; m331 = m331 + 1) 
        begin: inbit331
            assign data_11[m331 + b331*16 + a11*28*16] = data_11_array[a11][b331][m331];
        end
    endgenerate
    generate 
        localparam integer b332 = 24;
        for (m332 = 0; m332 < 16; m332 = m332 + 1) 
        begin: inbit332
            assign data_11[m332 + b332*16 + a11*28*16] = data_11_array[a11][b332][m332];
        end
    endgenerate
    generate 
        localparam integer b333 = 25;
        for (m333 = 0; m333 < 16; m333 = m333 + 1) 
        begin: inbit333
            assign data_11[m333 + b333*16 + a11*28*16] = data_11_array[a11][b333][m333];
        end
    endgenerate
    generate 
        localparam integer b334 = 26;
        for (m334 = 0; m334 < 16; m334 = m334 + 1) 
        begin: inbit334
            assign data_11[m334 + b334*16 + a11*28*16] = data_11_array[a11][b334][m334];
        end
    endgenerate
    generate 
        localparam integer b335 = 27;
        for (m335 = 0; m335 < 16; m335 = m335 + 1) 
        begin: inbit335
            assign data_11[m335 + b335*16 + a11*28*16] = data_11_array[a11][b335][m335];
        end
    endgenerate
    localparam integer a12 = 12;
    generate 
        localparam integer b336 = 0;
        for (m336 = 0; m336 < 16; m336 = m336 + 1) 
        begin: inbit336
            assign data_11[m336 + b336*16 + a12*28*16] = data_11_array[a12][b336][m336];
        end
    endgenerate
    generate 
        localparam integer b337 = 1;
        for (m337 = 0; m337 < 16; m337 = m337 + 1) 
        begin: inbit337
            assign data_11[m337 + b337*16 + a12*28*16] = data_11_array[a12][b337][m337];
        end
    endgenerate
    generate 
        localparam integer b338 = 2;
        for (m338 = 0; m338 < 16; m338 = m338 + 1) 
        begin: inbit338
            assign data_11[m338 + b338*16 + a12*28*16] = data_11_array[a12][b338][m338];
        end
    endgenerate
    generate 
        localparam integer b339 = 3;
        for (m339 = 0; m339 < 16; m339 = m339 + 1) 
        begin: inbit339
            assign data_11[m339 + b339*16 + a12*28*16] = data_11_array[a12][b339][m339];
        end
    endgenerate
    generate 
        localparam integer b340 = 4;
        for (m340 = 0; m340 < 16; m340 = m340 + 1) 
        begin: inbit340
            assign data_11[m340 + b340*16 + a12*28*16] = data_11_array[a12][b340][m340];
        end
    endgenerate
    generate 
        localparam integer b341 = 5;
        for (m341 = 0; m341 < 16; m341 = m341 + 1) 
        begin: inbit341
            assign data_11[m341 + b341*16 + a12*28*16] = data_11_array[a12][b341][m341];
        end
    endgenerate
    generate 
        localparam integer b342 = 6;
        for (m342 = 0; m342 < 16; m342 = m342 + 1) 
        begin: inbit342
            assign data_11[m342 + b342*16 + a12*28*16] = data_11_array[a12][b342][m342];
        end
    endgenerate
    generate 
        localparam integer b343 = 7;
        for (m343 = 0; m343 < 16; m343 = m343 + 1) 
        begin: inbit343
            assign data_11[m343 + b343*16 + a12*28*16] = data_11_array[a12][b343][m343];
        end
    endgenerate
    generate 
        localparam integer b344 = 8;
        for (m344 = 0; m344 < 16; m344 = m344 + 1) 
        begin: inbit344
            assign data_11[m344 + b344*16 + a12*28*16] = data_11_array[a12][b344][m344];
        end
    endgenerate
    generate 
        localparam integer b345 = 9;
        for (m345 = 0; m345 < 16; m345 = m345 + 1) 
        begin: inbit345
            assign data_11[m345 + b345*16 + a12*28*16] = data_11_array[a12][b345][m345];
        end
    endgenerate
    generate 
        localparam integer b346 = 10;
        for (m346 = 0; m346 < 16; m346 = m346 + 1) 
        begin: inbit346
            assign data_11[m346 + b346*16 + a12*28*16] = data_11_array[a12][b346][m346];
        end
    endgenerate
    generate 
        localparam integer b347 = 11;
        for (m347 = 0; m347 < 16; m347 = m347 + 1) 
        begin: inbit347
            assign data_11[m347 + b347*16 + a12*28*16] = data_11_array[a12][b347][m347];
        end
    endgenerate
    generate 
        localparam integer b348 = 12;
        for (m348 = 0; m348 < 16; m348 = m348 + 1) 
        begin: inbit348
            assign data_11[m348 + b348*16 + a12*28*16] = data_11_array[a12][b348][m348];
        end
    endgenerate
    generate 
        localparam integer b349 = 13;
        for (m349 = 0; m349 < 16; m349 = m349 + 1) 
        begin: inbit349
            assign data_11[m349 + b349*16 + a12*28*16] = data_11_array[a12][b349][m349];
        end
    endgenerate
    generate 
        localparam integer b350 = 14;
        for (m350 = 0; m350 < 16; m350 = m350 + 1) 
        begin: inbit350
            assign data_11[m350 + b350*16 + a12*28*16] = data_11_array[a12][b350][m350];
        end
    endgenerate
    generate 
        localparam integer b351 = 15;
        for (m351 = 0; m351 < 16; m351 = m351 + 1) 
        begin: inbit351
            assign data_11[m351 + b351*16 + a12*28*16] = data_11_array[a12][b351][m351];
        end
    endgenerate
    generate 
        localparam integer b352 = 16;
        for (m352 = 0; m352 < 16; m352 = m352 + 1) 
        begin: inbit352
            assign data_11[m352 + b352*16 + a12*28*16] = data_11_array[a12][b352][m352];
        end
    endgenerate
    generate 
        localparam integer b353 = 17;
        for (m353 = 0; m353 < 16; m353 = m353 + 1) 
        begin: inbit353
            assign data_11[m353 + b353*16 + a12*28*16] = data_11_array[a12][b353][m353];
        end
    endgenerate
    generate 
        localparam integer b354 = 18;
        for (m354 = 0; m354 < 16; m354 = m354 + 1) 
        begin: inbit354
            assign data_11[m354 + b354*16 + a12*28*16] = data_11_array[a12][b354][m354];
        end
    endgenerate
    generate 
        localparam integer b355 = 19;
        for (m355 = 0; m355 < 16; m355 = m355 + 1) 
        begin: inbit355
            assign data_11[m355 + b355*16 + a12*28*16] = data_11_array[a12][b355][m355];
        end
    endgenerate
    generate 
        localparam integer b356 = 20;
        for (m356 = 0; m356 < 16; m356 = m356 + 1) 
        begin: inbit356
            assign data_11[m356 + b356*16 + a12*28*16] = data_11_array[a12][b356][m356];
        end
    endgenerate
    generate 
        localparam integer b357 = 21;
        for (m357 = 0; m357 < 16; m357 = m357 + 1) 
        begin: inbit357
            assign data_11[m357 + b357*16 + a12*28*16] = data_11_array[a12][b357][m357];
        end
    endgenerate
    generate 
        localparam integer b358 = 22;
        for (m358 = 0; m358 < 16; m358 = m358 + 1) 
        begin: inbit358
            assign data_11[m358 + b358*16 + a12*28*16] = data_11_array[a12][b358][m358];
        end
    endgenerate
    generate 
        localparam integer b359 = 23;
        for (m359 = 0; m359 < 16; m359 = m359 + 1) 
        begin: inbit359
            assign data_11[m359 + b359*16 + a12*28*16] = data_11_array[a12][b359][m359];
        end
    endgenerate
    generate 
        localparam integer b360 = 24;
        for (m360 = 0; m360 < 16; m360 = m360 + 1) 
        begin: inbit360
            assign data_11[m360 + b360*16 + a12*28*16] = data_11_array[a12][b360][m360];
        end
    endgenerate
    generate 
        localparam integer b361 = 25;
        for (m361 = 0; m361 < 16; m361 = m361 + 1) 
        begin: inbit361
            assign data_11[m361 + b361*16 + a12*28*16] = data_11_array[a12][b361][m361];
        end
    endgenerate
    generate 
        localparam integer b362 = 26;
        for (m362 = 0; m362 < 16; m362 = m362 + 1) 
        begin: inbit362
            assign data_11[m362 + b362*16 + a12*28*16] = data_11_array[a12][b362][m362];
        end
    endgenerate
    generate 
        localparam integer b363 = 27;
        for (m363 = 0; m363 < 16; m363 = m363 + 1) 
        begin: inbit363
            assign data_11[m363 + b363*16 + a12*28*16] = data_11_array[a12][b363][m363];
        end
    endgenerate
    localparam integer a13 = 13;
    generate 
        localparam integer b364 = 0;
        for (m364 = 0; m364 < 16; m364 = m364 + 1) 
        begin: inbit364
            assign data_11[m364 + b364*16 + a13*28*16] = data_11_array[a13][b364][m364];
        end
    endgenerate
    generate 
        localparam integer b365 = 1;
        for (m365 = 0; m365 < 16; m365 = m365 + 1) 
        begin: inbit365
            assign data_11[m365 + b365*16 + a13*28*16] = data_11_array[a13][b365][m365];
        end
    endgenerate
    generate 
        localparam integer b366 = 2;
        for (m366 = 0; m366 < 16; m366 = m366 + 1) 
        begin: inbit366
            assign data_11[m366 + b366*16 + a13*28*16] = data_11_array[a13][b366][m366];
        end
    endgenerate
    generate 
        localparam integer b367 = 3;
        for (m367 = 0; m367 < 16; m367 = m367 + 1) 
        begin: inbit367
            assign data_11[m367 + b367*16 + a13*28*16] = data_11_array[a13][b367][m367];
        end
    endgenerate
    generate 
        localparam integer b368 = 4;
        for (m368 = 0; m368 < 16; m368 = m368 + 1) 
        begin: inbit368
            assign data_11[m368 + b368*16 + a13*28*16] = data_11_array[a13][b368][m368];
        end
    endgenerate
    generate 
        localparam integer b369 = 5;
        for (m369 = 0; m369 < 16; m369 = m369 + 1) 
        begin: inbit369
            assign data_11[m369 + b369*16 + a13*28*16] = data_11_array[a13][b369][m369];
        end
    endgenerate
    generate 
        localparam integer b370 = 6;
        for (m370 = 0; m370 < 16; m370 = m370 + 1) 
        begin: inbit370
            assign data_11[m370 + b370*16 + a13*28*16] = data_11_array[a13][b370][m370];
        end
    endgenerate
    generate 
        localparam integer b371 = 7;
        for (m371 = 0; m371 < 16; m371 = m371 + 1) 
        begin: inbit371
            assign data_11[m371 + b371*16 + a13*28*16] = data_11_array[a13][b371][m371];
        end
    endgenerate
    generate 
        localparam integer b372 = 8;
        for (m372 = 0; m372 < 16; m372 = m372 + 1) 
        begin: inbit372
            assign data_11[m372 + b372*16 + a13*28*16] = data_11_array[a13][b372][m372];
        end
    endgenerate
    generate 
        localparam integer b373 = 9;
        for (m373 = 0; m373 < 16; m373 = m373 + 1) 
        begin: inbit373
            assign data_11[m373 + b373*16 + a13*28*16] = data_11_array[a13][b373][m373];
        end
    endgenerate
    generate 
        localparam integer b374 = 10;
        for (m374 = 0; m374 < 16; m374 = m374 + 1) 
        begin: inbit374
            assign data_11[m374 + b374*16 + a13*28*16] = data_11_array[a13][b374][m374];
        end
    endgenerate
    generate 
        localparam integer b375 = 11;
        for (m375 = 0; m375 < 16; m375 = m375 + 1) 
        begin: inbit375
            assign data_11[m375 + b375*16 + a13*28*16] = data_11_array[a13][b375][m375];
        end
    endgenerate
    generate 
        localparam integer b376 = 12;
        for (m376 = 0; m376 < 16; m376 = m376 + 1) 
        begin: inbit376
            assign data_11[m376 + b376*16 + a13*28*16] = data_11_array[a13][b376][m376];
        end
    endgenerate
    generate 
        localparam integer b377 = 13;
        for (m377 = 0; m377 < 16; m377 = m377 + 1) 
        begin: inbit377
            assign data_11[m377 + b377*16 + a13*28*16] = data_11_array[a13][b377][m377];
        end
    endgenerate
    generate 
        localparam integer b378 = 14;
        for (m378 = 0; m378 < 16; m378 = m378 + 1) 
        begin: inbit378
            assign data_11[m378 + b378*16 + a13*28*16] = data_11_array[a13][b378][m378];
        end
    endgenerate
    generate 
        localparam integer b379 = 15;
        for (m379 = 0; m379 < 16; m379 = m379 + 1) 
        begin: inbit379
            assign data_11[m379 + b379*16 + a13*28*16] = data_11_array[a13][b379][m379];
        end
    endgenerate
    generate 
        localparam integer b380 = 16;
        for (m380 = 0; m380 < 16; m380 = m380 + 1) 
        begin: inbit380
            assign data_11[m380 + b380*16 + a13*28*16] = data_11_array[a13][b380][m380];
        end
    endgenerate
    generate 
        localparam integer b381 = 17;
        for (m381 = 0; m381 < 16; m381 = m381 + 1) 
        begin: inbit381
            assign data_11[m381 + b381*16 + a13*28*16] = data_11_array[a13][b381][m381];
        end
    endgenerate
    generate 
        localparam integer b382 = 18;
        for (m382 = 0; m382 < 16; m382 = m382 + 1) 
        begin: inbit382
            assign data_11[m382 + b382*16 + a13*28*16] = data_11_array[a13][b382][m382];
        end
    endgenerate
    generate 
        localparam integer b383 = 19;
        for (m383 = 0; m383 < 16; m383 = m383 + 1) 
        begin: inbit383
            assign data_11[m383 + b383*16 + a13*28*16] = data_11_array[a13][b383][m383];
        end
    endgenerate
    generate 
        localparam integer b384 = 20;
        for (m384 = 0; m384 < 16; m384 = m384 + 1) 
        begin: inbit384
            assign data_11[m384 + b384*16 + a13*28*16] = data_11_array[a13][b384][m384];
        end
    endgenerate
    generate 
        localparam integer b385 = 21;
        for (m385 = 0; m385 < 16; m385 = m385 + 1) 
        begin: inbit385
            assign data_11[m385 + b385*16 + a13*28*16] = data_11_array[a13][b385][m385];
        end
    endgenerate
    generate 
        localparam integer b386 = 22;
        for (m386 = 0; m386 < 16; m386 = m386 + 1) 
        begin: inbit386
            assign data_11[m386 + b386*16 + a13*28*16] = data_11_array[a13][b386][m386];
        end
    endgenerate
    generate 
        localparam integer b387 = 23;
        for (m387 = 0; m387 < 16; m387 = m387 + 1) 
        begin: inbit387
            assign data_11[m387 + b387*16 + a13*28*16] = data_11_array[a13][b387][m387];
        end
    endgenerate
    generate 
        localparam integer b388 = 24;
        for (m388 = 0; m388 < 16; m388 = m388 + 1) 
        begin: inbit388
            assign data_11[m388 + b388*16 + a13*28*16] = data_11_array[a13][b388][m388];
        end
    endgenerate
    generate 
        localparam integer b389 = 25;
        for (m389 = 0; m389 < 16; m389 = m389 + 1) 
        begin: inbit389
            assign data_11[m389 + b389*16 + a13*28*16] = data_11_array[a13][b389][m389];
        end
    endgenerate
    generate 
        localparam integer b390 = 26;
        for (m390 = 0; m390 < 16; m390 = m390 + 1) 
        begin: inbit390
            assign data_11[m390 + b390*16 + a13*28*16] = data_11_array[a13][b390][m390];
        end
    endgenerate
    generate 
        localparam integer b391 = 27;
        for (m391 = 0; m391 < 16; m391 = m391 + 1) 
        begin: inbit391
            assign data_11[m391 + b391*16 + a13*28*16] = data_11_array[a13][b391][m391];
        end
    endgenerate
    localparam integer a14 = 14;
    generate 
        localparam integer b392 = 0;
        for (m392 = 0; m392 < 16; m392 = m392 + 1) 
        begin: inbit392
            assign data_11[m392 + b392*16 + a14*28*16] = data_11_array[a14][b392][m392];
        end
    endgenerate
    generate 
        localparam integer b393 = 1;
        for (m393 = 0; m393 < 16; m393 = m393 + 1) 
        begin: inbit393
            assign data_11[m393 + b393*16 + a14*28*16] = data_11_array[a14][b393][m393];
        end
    endgenerate
    generate 
        localparam integer b394 = 2;
        for (m394 = 0; m394 < 16; m394 = m394 + 1) 
        begin: inbit394
            assign data_11[m394 + b394*16 + a14*28*16] = data_11_array[a14][b394][m394];
        end
    endgenerate
    generate 
        localparam integer b395 = 3;
        for (m395 = 0; m395 < 16; m395 = m395 + 1) 
        begin: inbit395
            assign data_11[m395 + b395*16 + a14*28*16] = data_11_array[a14][b395][m395];
        end
    endgenerate
    generate 
        localparam integer b396 = 4;
        for (m396 = 0; m396 < 16; m396 = m396 + 1) 
        begin: inbit396
            assign data_11[m396 + b396*16 + a14*28*16] = data_11_array[a14][b396][m396];
        end
    endgenerate
    generate 
        localparam integer b397 = 5;
        for (m397 = 0; m397 < 16; m397 = m397 + 1) 
        begin: inbit397
            assign data_11[m397 + b397*16 + a14*28*16] = data_11_array[a14][b397][m397];
        end
    endgenerate
    generate 
        localparam integer b398 = 6;
        for (m398 = 0; m398 < 16; m398 = m398 + 1) 
        begin: inbit398
            assign data_11[m398 + b398*16 + a14*28*16] = data_11_array[a14][b398][m398];
        end
    endgenerate
    generate 
        localparam integer b399 = 7;
        for (m399 = 0; m399 < 16; m399 = m399 + 1) 
        begin: inbit399
            assign data_11[m399 + b399*16 + a14*28*16] = data_11_array[a14][b399][m399];
        end
    endgenerate
    generate 
        localparam integer b400 = 8;
        for (m400 = 0; m400 < 16; m400 = m400 + 1) 
        begin: inbit400
            assign data_11[m400 + b400*16 + a14*28*16] = data_11_array[a14][b400][m400];
        end
    endgenerate
    generate 
        localparam integer b401 = 9;
        for (m401 = 0; m401 < 16; m401 = m401 + 1) 
        begin: inbit401
            assign data_11[m401 + b401*16 + a14*28*16] = data_11_array[a14][b401][m401];
        end
    endgenerate
    generate 
        localparam integer b402 = 10;
        for (m402 = 0; m402 < 16; m402 = m402 + 1) 
        begin: inbit402
            assign data_11[m402 + b402*16 + a14*28*16] = data_11_array[a14][b402][m402];
        end
    endgenerate
    generate 
        localparam integer b403 = 11;
        for (m403 = 0; m403 < 16; m403 = m403 + 1) 
        begin: inbit403
            assign data_11[m403 + b403*16 + a14*28*16] = data_11_array[a14][b403][m403];
        end
    endgenerate
    generate 
        localparam integer b404 = 12;
        for (m404 = 0; m404 < 16; m404 = m404 + 1) 
        begin: inbit404
            assign data_11[m404 + b404*16 + a14*28*16] = data_11_array[a14][b404][m404];
        end
    endgenerate
    generate 
        localparam integer b405 = 13;
        for (m405 = 0; m405 < 16; m405 = m405 + 1) 
        begin: inbit405
            assign data_11[m405 + b405*16 + a14*28*16] = data_11_array[a14][b405][m405];
        end
    endgenerate
    generate 
        localparam integer b406 = 14;
        for (m406 = 0; m406 < 16; m406 = m406 + 1) 
        begin: inbit406
            assign data_11[m406 + b406*16 + a14*28*16] = data_11_array[a14][b406][m406];
        end
    endgenerate
    generate 
        localparam integer b407 = 15;
        for (m407 = 0; m407 < 16; m407 = m407 + 1) 
        begin: inbit407
            assign data_11[m407 + b407*16 + a14*28*16] = data_11_array[a14][b407][m407];
        end
    endgenerate
    generate 
        localparam integer b408 = 16;
        for (m408 = 0; m408 < 16; m408 = m408 + 1) 
        begin: inbit408
            assign data_11[m408 + b408*16 + a14*28*16] = data_11_array[a14][b408][m408];
        end
    endgenerate
    generate 
        localparam integer b409 = 17;
        for (m409 = 0; m409 < 16; m409 = m409 + 1) 
        begin: inbit409
            assign data_11[m409 + b409*16 + a14*28*16] = data_11_array[a14][b409][m409];
        end
    endgenerate
    generate 
        localparam integer b410 = 18;
        for (m410 = 0; m410 < 16; m410 = m410 + 1) 
        begin: inbit410
            assign data_11[m410 + b410*16 + a14*28*16] = data_11_array[a14][b410][m410];
        end
    endgenerate
    generate 
        localparam integer b411 = 19;
        for (m411 = 0; m411 < 16; m411 = m411 + 1) 
        begin: inbit411
            assign data_11[m411 + b411*16 + a14*28*16] = data_11_array[a14][b411][m411];
        end
    endgenerate
    generate 
        localparam integer b412 = 20;
        for (m412 = 0; m412 < 16; m412 = m412 + 1) 
        begin: inbit412
            assign data_11[m412 + b412*16 + a14*28*16] = data_11_array[a14][b412][m412];
        end
    endgenerate
    generate 
        localparam integer b413 = 21;
        for (m413 = 0; m413 < 16; m413 = m413 + 1) 
        begin: inbit413
            assign data_11[m413 + b413*16 + a14*28*16] = data_11_array[a14][b413][m413];
        end
    endgenerate
    generate 
        localparam integer b414 = 22;
        for (m414 = 0; m414 < 16; m414 = m414 + 1) 
        begin: inbit414
            assign data_11[m414 + b414*16 + a14*28*16] = data_11_array[a14][b414][m414];
        end
    endgenerate
    generate 
        localparam integer b415 = 23;
        for (m415 = 0; m415 < 16; m415 = m415 + 1) 
        begin: inbit415
            assign data_11[m415 + b415*16 + a14*28*16] = data_11_array[a14][b415][m415];
        end
    endgenerate
    generate 
        localparam integer b416 = 24;
        for (m416 = 0; m416 < 16; m416 = m416 + 1) 
        begin: inbit416
            assign data_11[m416 + b416*16 + a14*28*16] = data_11_array[a14][b416][m416];
        end
    endgenerate
    generate 
        localparam integer b417 = 25;
        for (m417 = 0; m417 < 16; m417 = m417 + 1) 
        begin: inbit417
            assign data_11[m417 + b417*16 + a14*28*16] = data_11_array[a14][b417][m417];
        end
    endgenerate
    generate 
        localparam integer b418 = 26;
        for (m418 = 0; m418 < 16; m418 = m418 + 1) 
        begin: inbit418
            assign data_11[m418 + b418*16 + a14*28*16] = data_11_array[a14][b418][m418];
        end
    endgenerate
    generate 
        localparam integer b419 = 27;
        for (m419 = 0; m419 < 16; m419 = m419 + 1) 
        begin: inbit419
            assign data_11[m419 + b419*16 + a14*28*16] = data_11_array[a14][b419][m419];
        end
    endgenerate
    localparam integer a15 = 15;
    generate 
        localparam integer b420 = 0;
        for (m420 = 0; m420 < 16; m420 = m420 + 1) 
        begin: inbit420
            assign data_11[m420 + b420*16 + a15*28*16] = data_11_array[a15][b420][m420];
        end
    endgenerate
    generate 
        localparam integer b421 = 1;
        for (m421 = 0; m421 < 16; m421 = m421 + 1) 
        begin: inbit421
            assign data_11[m421 + b421*16 + a15*28*16] = data_11_array[a15][b421][m421];
        end
    endgenerate
    generate 
        localparam integer b422 = 2;
        for (m422 = 0; m422 < 16; m422 = m422 + 1) 
        begin: inbit422
            assign data_11[m422 + b422*16 + a15*28*16] = data_11_array[a15][b422][m422];
        end
    endgenerate
    generate 
        localparam integer b423 = 3;
        for (m423 = 0; m423 < 16; m423 = m423 + 1) 
        begin: inbit423
            assign data_11[m423 + b423*16 + a15*28*16] = data_11_array[a15][b423][m423];
        end
    endgenerate
    generate 
        localparam integer b424 = 4;
        for (m424 = 0; m424 < 16; m424 = m424 + 1) 
        begin: inbit424
            assign data_11[m424 + b424*16 + a15*28*16] = data_11_array[a15][b424][m424];
        end
    endgenerate
    generate 
        localparam integer b425 = 5;
        for (m425 = 0; m425 < 16; m425 = m425 + 1) 
        begin: inbit425
            assign data_11[m425 + b425*16 + a15*28*16] = data_11_array[a15][b425][m425];
        end
    endgenerate
    generate 
        localparam integer b426 = 6;
        for (m426 = 0; m426 < 16; m426 = m426 + 1) 
        begin: inbit426
            assign data_11[m426 + b426*16 + a15*28*16] = data_11_array[a15][b426][m426];
        end
    endgenerate
    generate 
        localparam integer b427 = 7;
        for (m427 = 0; m427 < 16; m427 = m427 + 1) 
        begin: inbit427
            assign data_11[m427 + b427*16 + a15*28*16] = data_11_array[a15][b427][m427];
        end
    endgenerate
    generate 
        localparam integer b428 = 8;
        for (m428 = 0; m428 < 16; m428 = m428 + 1) 
        begin: inbit428
            assign data_11[m428 + b428*16 + a15*28*16] = data_11_array[a15][b428][m428];
        end
    endgenerate
    generate 
        localparam integer b429 = 9;
        for (m429 = 0; m429 < 16; m429 = m429 + 1) 
        begin: inbit429
            assign data_11[m429 + b429*16 + a15*28*16] = data_11_array[a15][b429][m429];
        end
    endgenerate
    generate 
        localparam integer b430 = 10;
        for (m430 = 0; m430 < 16; m430 = m430 + 1) 
        begin: inbit430
            assign data_11[m430 + b430*16 + a15*28*16] = data_11_array[a15][b430][m430];
        end
    endgenerate
    generate 
        localparam integer b431 = 11;
        for (m431 = 0; m431 < 16; m431 = m431 + 1) 
        begin: inbit431
            assign data_11[m431 + b431*16 + a15*28*16] = data_11_array[a15][b431][m431];
        end
    endgenerate
    generate 
        localparam integer b432 = 12;
        for (m432 = 0; m432 < 16; m432 = m432 + 1) 
        begin: inbit432
            assign data_11[m432 + b432*16 + a15*28*16] = data_11_array[a15][b432][m432];
        end
    endgenerate
    generate 
        localparam integer b433 = 13;
        for (m433 = 0; m433 < 16; m433 = m433 + 1) 
        begin: inbit433
            assign data_11[m433 + b433*16 + a15*28*16] = data_11_array[a15][b433][m433];
        end
    endgenerate
    generate 
        localparam integer b434 = 14;
        for (m434 = 0; m434 < 16; m434 = m434 + 1) 
        begin: inbit434
            assign data_11[m434 + b434*16 + a15*28*16] = data_11_array[a15][b434][m434];
        end
    endgenerate
    generate 
        localparam integer b435 = 15;
        for (m435 = 0; m435 < 16; m435 = m435 + 1) 
        begin: inbit435
            assign data_11[m435 + b435*16 + a15*28*16] = data_11_array[a15][b435][m435];
        end
    endgenerate
    generate 
        localparam integer b436 = 16;
        for (m436 = 0; m436 < 16; m436 = m436 + 1) 
        begin: inbit436
            assign data_11[m436 + b436*16 + a15*28*16] = data_11_array[a15][b436][m436];
        end
    endgenerate
    generate 
        localparam integer b437 = 17;
        for (m437 = 0; m437 < 16; m437 = m437 + 1) 
        begin: inbit437
            assign data_11[m437 + b437*16 + a15*28*16] = data_11_array[a15][b437][m437];
        end
    endgenerate
    generate 
        localparam integer b438 = 18;
        for (m438 = 0; m438 < 16; m438 = m438 + 1) 
        begin: inbit438
            assign data_11[m438 + b438*16 + a15*28*16] = data_11_array[a15][b438][m438];
        end
    endgenerate
    generate 
        localparam integer b439 = 19;
        for (m439 = 0; m439 < 16; m439 = m439 + 1) 
        begin: inbit439
            assign data_11[m439 + b439*16 + a15*28*16] = data_11_array[a15][b439][m439];
        end
    endgenerate
    generate 
        localparam integer b440 = 20;
        for (m440 = 0; m440 < 16; m440 = m440 + 1) 
        begin: inbit440
            assign data_11[m440 + b440*16 + a15*28*16] = data_11_array[a15][b440][m440];
        end
    endgenerate
    generate 
        localparam integer b441 = 21;
        for (m441 = 0; m441 < 16; m441 = m441 + 1) 
        begin: inbit441
            assign data_11[m441 + b441*16 + a15*28*16] = data_11_array[a15][b441][m441];
        end
    endgenerate
    generate 
        localparam integer b442 = 22;
        for (m442 = 0; m442 < 16; m442 = m442 + 1) 
        begin: inbit442
            assign data_11[m442 + b442*16 + a15*28*16] = data_11_array[a15][b442][m442];
        end
    endgenerate
    generate 
        localparam integer b443 = 23;
        for (m443 = 0; m443 < 16; m443 = m443 + 1) 
        begin: inbit443
            assign data_11[m443 + b443*16 + a15*28*16] = data_11_array[a15][b443][m443];
        end
    endgenerate
    generate 
        localparam integer b444 = 24;
        for (m444 = 0; m444 < 16; m444 = m444 + 1) 
        begin: inbit444
            assign data_11[m444 + b444*16 + a15*28*16] = data_11_array[a15][b444][m444];
        end
    endgenerate
    generate 
        localparam integer b445 = 25;
        for (m445 = 0; m445 < 16; m445 = m445 + 1) 
        begin: inbit445
            assign data_11[m445 + b445*16 + a15*28*16] = data_11_array[a15][b445][m445];
        end
    endgenerate
    generate 
        localparam integer b446 = 26;
        for (m446 = 0; m446 < 16; m446 = m446 + 1) 
        begin: inbit446
            assign data_11[m446 + b446*16 + a15*28*16] = data_11_array[a15][b446][m446];
        end
    endgenerate
    generate 
        localparam integer b447 = 27;
        for (m447 = 0; m447 < 16; m447 = m447 + 1) 
        begin: inbit447
            assign data_11[m447 + b447*16 + a15*28*16] = data_11_array[a15][b447][m447];
        end
    endgenerate
    localparam integer a16 = 16;
    generate 
        localparam integer b448 = 0;
        for (m448 = 0; m448 < 16; m448 = m448 + 1) 
        begin: inbit448
            assign data_11[m448 + b448*16 + a16*28*16] = data_11_array[a16][b448][m448];
        end
    endgenerate
    generate 
        localparam integer b449 = 1;
        for (m449 = 0; m449 < 16; m449 = m449 + 1) 
        begin: inbit449
            assign data_11[m449 + b449*16 + a16*28*16] = data_11_array[a16][b449][m449];
        end
    endgenerate
    generate 
        localparam integer b450 = 2;
        for (m450 = 0; m450 < 16; m450 = m450 + 1) 
        begin: inbit450
            assign data_11[m450 + b450*16 + a16*28*16] = data_11_array[a16][b450][m450];
        end
    endgenerate
    generate 
        localparam integer b451 = 3;
        for (m451 = 0; m451 < 16; m451 = m451 + 1) 
        begin: inbit451
            assign data_11[m451 + b451*16 + a16*28*16] = data_11_array[a16][b451][m451];
        end
    endgenerate
    generate 
        localparam integer b452 = 4;
        for (m452 = 0; m452 < 16; m452 = m452 + 1) 
        begin: inbit452
            assign data_11[m452 + b452*16 + a16*28*16] = data_11_array[a16][b452][m452];
        end
    endgenerate
    generate 
        localparam integer b453 = 5;
        for (m453 = 0; m453 < 16; m453 = m453 + 1) 
        begin: inbit453
            assign data_11[m453 + b453*16 + a16*28*16] = data_11_array[a16][b453][m453];
        end
    endgenerate
    generate 
        localparam integer b454 = 6;
        for (m454 = 0; m454 < 16; m454 = m454 + 1) 
        begin: inbit454
            assign data_11[m454 + b454*16 + a16*28*16] = data_11_array[a16][b454][m454];
        end
    endgenerate
    generate 
        localparam integer b455 = 7;
        for (m455 = 0; m455 < 16; m455 = m455 + 1) 
        begin: inbit455
            assign data_11[m455 + b455*16 + a16*28*16] = data_11_array[a16][b455][m455];
        end
    endgenerate
    generate 
        localparam integer b456 = 8;
        for (m456 = 0; m456 < 16; m456 = m456 + 1) 
        begin: inbit456
            assign data_11[m456 + b456*16 + a16*28*16] = data_11_array[a16][b456][m456];
        end
    endgenerate
    generate 
        localparam integer b457 = 9;
        for (m457 = 0; m457 < 16; m457 = m457 + 1) 
        begin: inbit457
            assign data_11[m457 + b457*16 + a16*28*16] = data_11_array[a16][b457][m457];
        end
    endgenerate
    generate 
        localparam integer b458 = 10;
        for (m458 = 0; m458 < 16; m458 = m458 + 1) 
        begin: inbit458
            assign data_11[m458 + b458*16 + a16*28*16] = data_11_array[a16][b458][m458];
        end
    endgenerate
    generate 
        localparam integer b459 = 11;
        for (m459 = 0; m459 < 16; m459 = m459 + 1) 
        begin: inbit459
            assign data_11[m459 + b459*16 + a16*28*16] = data_11_array[a16][b459][m459];
        end
    endgenerate
    generate 
        localparam integer b460 = 12;
        for (m460 = 0; m460 < 16; m460 = m460 + 1) 
        begin: inbit460
            assign data_11[m460 + b460*16 + a16*28*16] = data_11_array[a16][b460][m460];
        end
    endgenerate
    generate 
        localparam integer b461 = 13;
        for (m461 = 0; m461 < 16; m461 = m461 + 1) 
        begin: inbit461
            assign data_11[m461 + b461*16 + a16*28*16] = data_11_array[a16][b461][m461];
        end
    endgenerate
    generate 
        localparam integer b462 = 14;
        for (m462 = 0; m462 < 16; m462 = m462 + 1) 
        begin: inbit462
            assign data_11[m462 + b462*16 + a16*28*16] = data_11_array[a16][b462][m462];
        end
    endgenerate
    generate 
        localparam integer b463 = 15;
        for (m463 = 0; m463 < 16; m463 = m463 + 1) 
        begin: inbit463
            assign data_11[m463 + b463*16 + a16*28*16] = data_11_array[a16][b463][m463];
        end
    endgenerate
    generate 
        localparam integer b464 = 16;
        for (m464 = 0; m464 < 16; m464 = m464 + 1) 
        begin: inbit464
            assign data_11[m464 + b464*16 + a16*28*16] = data_11_array[a16][b464][m464];
        end
    endgenerate
    generate 
        localparam integer b465 = 17;
        for (m465 = 0; m465 < 16; m465 = m465 + 1) 
        begin: inbit465
            assign data_11[m465 + b465*16 + a16*28*16] = data_11_array[a16][b465][m465];
        end
    endgenerate
    generate 
        localparam integer b466 = 18;
        for (m466 = 0; m466 < 16; m466 = m466 + 1) 
        begin: inbit466
            assign data_11[m466 + b466*16 + a16*28*16] = data_11_array[a16][b466][m466];
        end
    endgenerate
    generate 
        localparam integer b467 = 19;
        for (m467 = 0; m467 < 16; m467 = m467 + 1) 
        begin: inbit467
            assign data_11[m467 + b467*16 + a16*28*16] = data_11_array[a16][b467][m467];
        end
    endgenerate
    generate 
        localparam integer b468 = 20;
        for (m468 = 0; m468 < 16; m468 = m468 + 1) 
        begin: inbit468
            assign data_11[m468 + b468*16 + a16*28*16] = data_11_array[a16][b468][m468];
        end
    endgenerate
    generate 
        localparam integer b469 = 21;
        for (m469 = 0; m469 < 16; m469 = m469 + 1) 
        begin: inbit469
            assign data_11[m469 + b469*16 + a16*28*16] = data_11_array[a16][b469][m469];
        end
    endgenerate
    generate 
        localparam integer b470 = 22;
        for (m470 = 0; m470 < 16; m470 = m470 + 1) 
        begin: inbit470
            assign data_11[m470 + b470*16 + a16*28*16] = data_11_array[a16][b470][m470];
        end
    endgenerate
    generate 
        localparam integer b471 = 23;
        for (m471 = 0; m471 < 16; m471 = m471 + 1) 
        begin: inbit471
            assign data_11[m471 + b471*16 + a16*28*16] = data_11_array[a16][b471][m471];
        end
    endgenerate
    generate 
        localparam integer b472 = 24;
        for (m472 = 0; m472 < 16; m472 = m472 + 1) 
        begin: inbit472
            assign data_11[m472 + b472*16 + a16*28*16] = data_11_array[a16][b472][m472];
        end
    endgenerate
    generate 
        localparam integer b473 = 25;
        for (m473 = 0; m473 < 16; m473 = m473 + 1) 
        begin: inbit473
            assign data_11[m473 + b473*16 + a16*28*16] = data_11_array[a16][b473][m473];
        end
    endgenerate
    generate 
        localparam integer b474 = 26;
        for (m474 = 0; m474 < 16; m474 = m474 + 1) 
        begin: inbit474
            assign data_11[m474 + b474*16 + a16*28*16] = data_11_array[a16][b474][m474];
        end
    endgenerate
    generate 
        localparam integer b475 = 27;
        for (m475 = 0; m475 < 16; m475 = m475 + 1) 
        begin: inbit475
            assign data_11[m475 + b475*16 + a16*28*16] = data_11_array[a16][b475][m475];
        end
    endgenerate
    localparam integer a17 = 17;
    generate 
        localparam integer b476 = 0;
        for (m476 = 0; m476 < 16; m476 = m476 + 1) 
        begin: inbit476
            assign data_11[m476 + b476*16 + a17*28*16] = data_11_array[a17][b476][m476];
        end
    endgenerate
    generate 
        localparam integer b477 = 1;
        for (m477 = 0; m477 < 16; m477 = m477 + 1) 
        begin: inbit477
            assign data_11[m477 + b477*16 + a17*28*16] = data_11_array[a17][b477][m477];
        end
    endgenerate
    generate 
        localparam integer b478 = 2;
        for (m478 = 0; m478 < 16; m478 = m478 + 1) 
        begin: inbit478
            assign data_11[m478 + b478*16 + a17*28*16] = data_11_array[a17][b478][m478];
        end
    endgenerate
    generate 
        localparam integer b479 = 3;
        for (m479 = 0; m479 < 16; m479 = m479 + 1) 
        begin: inbit479
            assign data_11[m479 + b479*16 + a17*28*16] = data_11_array[a17][b479][m479];
        end
    endgenerate
    generate 
        localparam integer b480 = 4;
        for (m480 = 0; m480 < 16; m480 = m480 + 1) 
        begin: inbit480
            assign data_11[m480 + b480*16 + a17*28*16] = data_11_array[a17][b480][m480];
        end
    endgenerate
    generate 
        localparam integer b481 = 5;
        for (m481 = 0; m481 < 16; m481 = m481 + 1) 
        begin: inbit481
            assign data_11[m481 + b481*16 + a17*28*16] = data_11_array[a17][b481][m481];
        end
    endgenerate
    generate 
        localparam integer b482 = 6;
        for (m482 = 0; m482 < 16; m482 = m482 + 1) 
        begin: inbit482
            assign data_11[m482 + b482*16 + a17*28*16] = data_11_array[a17][b482][m482];
        end
    endgenerate
    generate 
        localparam integer b483 = 7;
        for (m483 = 0; m483 < 16; m483 = m483 + 1) 
        begin: inbit483
            assign data_11[m483 + b483*16 + a17*28*16] = data_11_array[a17][b483][m483];
        end
    endgenerate
    generate 
        localparam integer b484 = 8;
        for (m484 = 0; m484 < 16; m484 = m484 + 1) 
        begin: inbit484
            assign data_11[m484 + b484*16 + a17*28*16] = data_11_array[a17][b484][m484];
        end
    endgenerate
    generate 
        localparam integer b485 = 9;
        for (m485 = 0; m485 < 16; m485 = m485 + 1) 
        begin: inbit485
            assign data_11[m485 + b485*16 + a17*28*16] = data_11_array[a17][b485][m485];
        end
    endgenerate
    generate 
        localparam integer b486 = 10;
        for (m486 = 0; m486 < 16; m486 = m486 + 1) 
        begin: inbit486
            assign data_11[m486 + b486*16 + a17*28*16] = data_11_array[a17][b486][m486];
        end
    endgenerate
    generate 
        localparam integer b487 = 11;
        for (m487 = 0; m487 < 16; m487 = m487 + 1) 
        begin: inbit487
            assign data_11[m487 + b487*16 + a17*28*16] = data_11_array[a17][b487][m487];
        end
    endgenerate
    generate 
        localparam integer b488 = 12;
        for (m488 = 0; m488 < 16; m488 = m488 + 1) 
        begin: inbit488
            assign data_11[m488 + b488*16 + a17*28*16] = data_11_array[a17][b488][m488];
        end
    endgenerate
    generate 
        localparam integer b489 = 13;
        for (m489 = 0; m489 < 16; m489 = m489 + 1) 
        begin: inbit489
            assign data_11[m489 + b489*16 + a17*28*16] = data_11_array[a17][b489][m489];
        end
    endgenerate
    generate 
        localparam integer b490 = 14;
        for (m490 = 0; m490 < 16; m490 = m490 + 1) 
        begin: inbit490
            assign data_11[m490 + b490*16 + a17*28*16] = data_11_array[a17][b490][m490];
        end
    endgenerate
    generate 
        localparam integer b491 = 15;
        for (m491 = 0; m491 < 16; m491 = m491 + 1) 
        begin: inbit491
            assign data_11[m491 + b491*16 + a17*28*16] = data_11_array[a17][b491][m491];
        end
    endgenerate
    generate 
        localparam integer b492 = 16;
        for (m492 = 0; m492 < 16; m492 = m492 + 1) 
        begin: inbit492
            assign data_11[m492 + b492*16 + a17*28*16] = data_11_array[a17][b492][m492];
        end
    endgenerate
    generate 
        localparam integer b493 = 17;
        for (m493 = 0; m493 < 16; m493 = m493 + 1) 
        begin: inbit493
            assign data_11[m493 + b493*16 + a17*28*16] = data_11_array[a17][b493][m493];
        end
    endgenerate
    generate 
        localparam integer b494 = 18;
        for (m494 = 0; m494 < 16; m494 = m494 + 1) 
        begin: inbit494
            assign data_11[m494 + b494*16 + a17*28*16] = data_11_array[a17][b494][m494];
        end
    endgenerate
    generate 
        localparam integer b495 = 19;
        for (m495 = 0; m495 < 16; m495 = m495 + 1) 
        begin: inbit495
            assign data_11[m495 + b495*16 + a17*28*16] = data_11_array[a17][b495][m495];
        end
    endgenerate
    generate 
        localparam integer b496 = 20;
        for (m496 = 0; m496 < 16; m496 = m496 + 1) 
        begin: inbit496
            assign data_11[m496 + b496*16 + a17*28*16] = data_11_array[a17][b496][m496];
        end
    endgenerate
    generate 
        localparam integer b497 = 21;
        for (m497 = 0; m497 < 16; m497 = m497 + 1) 
        begin: inbit497
            assign data_11[m497 + b497*16 + a17*28*16] = data_11_array[a17][b497][m497];
        end
    endgenerate
    generate 
        localparam integer b498 = 22;
        for (m498 = 0; m498 < 16; m498 = m498 + 1) 
        begin: inbit498
            assign data_11[m498 + b498*16 + a17*28*16] = data_11_array[a17][b498][m498];
        end
    endgenerate
    generate 
        localparam integer b499 = 23;
        for (m499 = 0; m499 < 16; m499 = m499 + 1) 
        begin: inbit499
            assign data_11[m499 + b499*16 + a17*28*16] = data_11_array[a17][b499][m499];
        end
    endgenerate
    generate 
        localparam integer b500 = 24;
        for (m500 = 0; m500 < 16; m500 = m500 + 1) 
        begin: inbit500
            assign data_11[m500 + b500*16 + a17*28*16] = data_11_array[a17][b500][m500];
        end
    endgenerate
    generate 
        localparam integer b501 = 25;
        for (m501 = 0; m501 < 16; m501 = m501 + 1) 
        begin: inbit501
            assign data_11[m501 + b501*16 + a17*28*16] = data_11_array[a17][b501][m501];
        end
    endgenerate
    generate 
        localparam integer b502 = 26;
        for (m502 = 0; m502 < 16; m502 = m502 + 1) 
        begin: inbit502
            assign data_11[m502 + b502*16 + a17*28*16] = data_11_array[a17][b502][m502];
        end
    endgenerate
    generate 
        localparam integer b503 = 27;
        for (m503 = 0; m503 < 16; m503 = m503 + 1) 
        begin: inbit503
            assign data_11[m503 + b503*16 + a17*28*16] = data_11_array[a17][b503][m503];
        end
    endgenerate
    localparam integer a18 = 18;
    generate 
        localparam integer b504 = 0;
        for (m504 = 0; m504 < 16; m504 = m504 + 1) 
        begin: inbit504
            assign data_11[m504 + b504*16 + a18*28*16] = data_11_array[a18][b504][m504];
        end
    endgenerate
    generate 
        localparam integer b505 = 1;
        for (m505 = 0; m505 < 16; m505 = m505 + 1) 
        begin: inbit505
            assign data_11[m505 + b505*16 + a18*28*16] = data_11_array[a18][b505][m505];
        end
    endgenerate
    generate 
        localparam integer b506 = 2;
        for (m506 = 0; m506 < 16; m506 = m506 + 1) 
        begin: inbit506
            assign data_11[m506 + b506*16 + a18*28*16] = data_11_array[a18][b506][m506];
        end
    endgenerate
    generate 
        localparam integer b507 = 3;
        for (m507 = 0; m507 < 16; m507 = m507 + 1) 
        begin: inbit507
            assign data_11[m507 + b507*16 + a18*28*16] = data_11_array[a18][b507][m507];
        end
    endgenerate
    generate 
        localparam integer b508 = 4;
        for (m508 = 0; m508 < 16; m508 = m508 + 1) 
        begin: inbit508
            assign data_11[m508 + b508*16 + a18*28*16] = data_11_array[a18][b508][m508];
        end
    endgenerate
    generate 
        localparam integer b509 = 5;
        for (m509 = 0; m509 < 16; m509 = m509 + 1) 
        begin: inbit509
            assign data_11[m509 + b509*16 + a18*28*16] = data_11_array[a18][b509][m509];
        end
    endgenerate
    generate 
        localparam integer b510 = 6;
        for (m510 = 0; m510 < 16; m510 = m510 + 1) 
        begin: inbit510
            assign data_11[m510 + b510*16 + a18*28*16] = data_11_array[a18][b510][m510];
        end
    endgenerate
    generate 
        localparam integer b511 = 7;
        for (m511 = 0; m511 < 16; m511 = m511 + 1) 
        begin: inbit511
            assign data_11[m511 + b511*16 + a18*28*16] = data_11_array[a18][b511][m511];
        end
    endgenerate
    generate 
        localparam integer b512 = 8;
        for (m512 = 0; m512 < 16; m512 = m512 + 1) 
        begin: inbit512
            assign data_11[m512 + b512*16 + a18*28*16] = data_11_array[a18][b512][m512];
        end
    endgenerate
    generate 
        localparam integer b513 = 9;
        for (m513 = 0; m513 < 16; m513 = m513 + 1) 
        begin: inbit513
            assign data_11[m513 + b513*16 + a18*28*16] = data_11_array[a18][b513][m513];
        end
    endgenerate
    generate 
        localparam integer b514 = 10;
        for (m514 = 0; m514 < 16; m514 = m514 + 1) 
        begin: inbit514
            assign data_11[m514 + b514*16 + a18*28*16] = data_11_array[a18][b514][m514];
        end
    endgenerate
    generate 
        localparam integer b515 = 11;
        for (m515 = 0; m515 < 16; m515 = m515 + 1) 
        begin: inbit515
            assign data_11[m515 + b515*16 + a18*28*16] = data_11_array[a18][b515][m515];
        end
    endgenerate
    generate 
        localparam integer b516 = 12;
        for (m516 = 0; m516 < 16; m516 = m516 + 1) 
        begin: inbit516
            assign data_11[m516 + b516*16 + a18*28*16] = data_11_array[a18][b516][m516];
        end
    endgenerate
    generate 
        localparam integer b517 = 13;
        for (m517 = 0; m517 < 16; m517 = m517 + 1) 
        begin: inbit517
            assign data_11[m517 + b517*16 + a18*28*16] = data_11_array[a18][b517][m517];
        end
    endgenerate
    generate 
        localparam integer b518 = 14;
        for (m518 = 0; m518 < 16; m518 = m518 + 1) 
        begin: inbit518
            assign data_11[m518 + b518*16 + a18*28*16] = data_11_array[a18][b518][m518];
        end
    endgenerate
    generate 
        localparam integer b519 = 15;
        for (m519 = 0; m519 < 16; m519 = m519 + 1) 
        begin: inbit519
            assign data_11[m519 + b519*16 + a18*28*16] = data_11_array[a18][b519][m519];
        end
    endgenerate
    generate 
        localparam integer b520 = 16;
        for (m520 = 0; m520 < 16; m520 = m520 + 1) 
        begin: inbit520
            assign data_11[m520 + b520*16 + a18*28*16] = data_11_array[a18][b520][m520];
        end
    endgenerate
    generate 
        localparam integer b521 = 17;
        for (m521 = 0; m521 < 16; m521 = m521 + 1) 
        begin: inbit521
            assign data_11[m521 + b521*16 + a18*28*16] = data_11_array[a18][b521][m521];
        end
    endgenerate
    generate 
        localparam integer b522 = 18;
        for (m522 = 0; m522 < 16; m522 = m522 + 1) 
        begin: inbit522
            assign data_11[m522 + b522*16 + a18*28*16] = data_11_array[a18][b522][m522];
        end
    endgenerate
    generate 
        localparam integer b523 = 19;
        for (m523 = 0; m523 < 16; m523 = m523 + 1) 
        begin: inbit523
            assign data_11[m523 + b523*16 + a18*28*16] = data_11_array[a18][b523][m523];
        end
    endgenerate
    generate 
        localparam integer b524 = 20;
        for (m524 = 0; m524 < 16; m524 = m524 + 1) 
        begin: inbit524
            assign data_11[m524 + b524*16 + a18*28*16] = data_11_array[a18][b524][m524];
        end
    endgenerate
    generate 
        localparam integer b525 = 21;
        for (m525 = 0; m525 < 16; m525 = m525 + 1) 
        begin: inbit525
            assign data_11[m525 + b525*16 + a18*28*16] = data_11_array[a18][b525][m525];
        end
    endgenerate
    generate 
        localparam integer b526 = 22;
        for (m526 = 0; m526 < 16; m526 = m526 + 1) 
        begin: inbit526
            assign data_11[m526 + b526*16 + a18*28*16] = data_11_array[a18][b526][m526];
        end
    endgenerate
    generate 
        localparam integer b527 = 23;
        for (m527 = 0; m527 < 16; m527 = m527 + 1) 
        begin: inbit527
            assign data_11[m527 + b527*16 + a18*28*16] = data_11_array[a18][b527][m527];
        end
    endgenerate
    generate 
        localparam integer b528 = 24;
        for (m528 = 0; m528 < 16; m528 = m528 + 1) 
        begin: inbit528
            assign data_11[m528 + b528*16 + a18*28*16] = data_11_array[a18][b528][m528];
        end
    endgenerate
    generate 
        localparam integer b529 = 25;
        for (m529 = 0; m529 < 16; m529 = m529 + 1) 
        begin: inbit529
            assign data_11[m529 + b529*16 + a18*28*16] = data_11_array[a18][b529][m529];
        end
    endgenerate
    generate 
        localparam integer b530 = 26;
        for (m530 = 0; m530 < 16; m530 = m530 + 1) 
        begin: inbit530
            assign data_11[m530 + b530*16 + a18*28*16] = data_11_array[a18][b530][m530];
        end
    endgenerate
    generate 
        localparam integer b531 = 27;
        for (m531 = 0; m531 < 16; m531 = m531 + 1) 
        begin: inbit531
            assign data_11[m531 + b531*16 + a18*28*16] = data_11_array[a18][b531][m531];
        end
    endgenerate
    localparam integer a19 = 19;
    generate 
        localparam integer b532 = 0;
        for (m532 = 0; m532 < 16; m532 = m532 + 1) 
        begin: inbit532
            assign data_11[m532 + b532*16 + a19*28*16] = data_11_array[a19][b532][m532];
        end
    endgenerate
    generate 
        localparam integer b533 = 1;
        for (m533 = 0; m533 < 16; m533 = m533 + 1) 
        begin: inbit533
            assign data_11[m533 + b533*16 + a19*28*16] = data_11_array[a19][b533][m533];
        end
    endgenerate
    generate 
        localparam integer b534 = 2;
        for (m534 = 0; m534 < 16; m534 = m534 + 1) 
        begin: inbit534
            assign data_11[m534 + b534*16 + a19*28*16] = data_11_array[a19][b534][m534];
        end
    endgenerate
    generate 
        localparam integer b535 = 3;
        for (m535 = 0; m535 < 16; m535 = m535 + 1) 
        begin: inbit535
            assign data_11[m535 + b535*16 + a19*28*16] = data_11_array[a19][b535][m535];
        end
    endgenerate
    generate 
        localparam integer b536 = 4;
        for (m536 = 0; m536 < 16; m536 = m536 + 1) 
        begin: inbit536
            assign data_11[m536 + b536*16 + a19*28*16] = data_11_array[a19][b536][m536];
        end
    endgenerate
    generate 
        localparam integer b537 = 5;
        for (m537 = 0; m537 < 16; m537 = m537 + 1) 
        begin: inbit537
            assign data_11[m537 + b537*16 + a19*28*16] = data_11_array[a19][b537][m537];
        end
    endgenerate
    generate 
        localparam integer b538 = 6;
        for (m538 = 0; m538 < 16; m538 = m538 + 1) 
        begin: inbit538
            assign data_11[m538 + b538*16 + a19*28*16] = data_11_array[a19][b538][m538];
        end
    endgenerate
    generate 
        localparam integer b539 = 7;
        for (m539 = 0; m539 < 16; m539 = m539 + 1) 
        begin: inbit539
            assign data_11[m539 + b539*16 + a19*28*16] = data_11_array[a19][b539][m539];
        end
    endgenerate
    generate 
        localparam integer b540 = 8;
        for (m540 = 0; m540 < 16; m540 = m540 + 1) 
        begin: inbit540
            assign data_11[m540 + b540*16 + a19*28*16] = data_11_array[a19][b540][m540];
        end
    endgenerate
    generate 
        localparam integer b541 = 9;
        for (m541 = 0; m541 < 16; m541 = m541 + 1) 
        begin: inbit541
            assign data_11[m541 + b541*16 + a19*28*16] = data_11_array[a19][b541][m541];
        end
    endgenerate
    generate 
        localparam integer b542 = 10;
        for (m542 = 0; m542 < 16; m542 = m542 + 1) 
        begin: inbit542
            assign data_11[m542 + b542*16 + a19*28*16] = data_11_array[a19][b542][m542];
        end
    endgenerate
    generate 
        localparam integer b543 = 11;
        for (m543 = 0; m543 < 16; m543 = m543 + 1) 
        begin: inbit543
            assign data_11[m543 + b543*16 + a19*28*16] = data_11_array[a19][b543][m543];
        end
    endgenerate
    generate 
        localparam integer b544 = 12;
        for (m544 = 0; m544 < 16; m544 = m544 + 1) 
        begin: inbit544
            assign data_11[m544 + b544*16 + a19*28*16] = data_11_array[a19][b544][m544];
        end
    endgenerate
    generate 
        localparam integer b545 = 13;
        for (m545 = 0; m545 < 16; m545 = m545 + 1) 
        begin: inbit545
            assign data_11[m545 + b545*16 + a19*28*16] = data_11_array[a19][b545][m545];
        end
    endgenerate
    generate 
        localparam integer b546 = 14;
        for (m546 = 0; m546 < 16; m546 = m546 + 1) 
        begin: inbit546
            assign data_11[m546 + b546*16 + a19*28*16] = data_11_array[a19][b546][m546];
        end
    endgenerate
    generate 
        localparam integer b547 = 15;
        for (m547 = 0; m547 < 16; m547 = m547 + 1) 
        begin: inbit547
            assign data_11[m547 + b547*16 + a19*28*16] = data_11_array[a19][b547][m547];
        end
    endgenerate
    generate 
        localparam integer b548 = 16;
        for (m548 = 0; m548 < 16; m548 = m548 + 1) 
        begin: inbit548
            assign data_11[m548 + b548*16 + a19*28*16] = data_11_array[a19][b548][m548];
        end
    endgenerate
    generate 
        localparam integer b549 = 17;
        for (m549 = 0; m549 < 16; m549 = m549 + 1) 
        begin: inbit549
            assign data_11[m549 + b549*16 + a19*28*16] = data_11_array[a19][b549][m549];
        end
    endgenerate
    generate 
        localparam integer b550 = 18;
        for (m550 = 0; m550 < 16; m550 = m550 + 1) 
        begin: inbit550
            assign data_11[m550 + b550*16 + a19*28*16] = data_11_array[a19][b550][m550];
        end
    endgenerate
    generate 
        localparam integer b551 = 19;
        for (m551 = 0; m551 < 16; m551 = m551 + 1) 
        begin: inbit551
            assign data_11[m551 + b551*16 + a19*28*16] = data_11_array[a19][b551][m551];
        end
    endgenerate
    generate 
        localparam integer b552 = 20;
        for (m552 = 0; m552 < 16; m552 = m552 + 1) 
        begin: inbit552
            assign data_11[m552 + b552*16 + a19*28*16] = data_11_array[a19][b552][m552];
        end
    endgenerate
    generate 
        localparam integer b553 = 21;
        for (m553 = 0; m553 < 16; m553 = m553 + 1) 
        begin: inbit553
            assign data_11[m553 + b553*16 + a19*28*16] = data_11_array[a19][b553][m553];
        end
    endgenerate
    generate 
        localparam integer b554 = 22;
        for (m554 = 0; m554 < 16; m554 = m554 + 1) 
        begin: inbit554
            assign data_11[m554 + b554*16 + a19*28*16] = data_11_array[a19][b554][m554];
        end
    endgenerate
    generate 
        localparam integer b555 = 23;
        for (m555 = 0; m555 < 16; m555 = m555 + 1) 
        begin: inbit555
            assign data_11[m555 + b555*16 + a19*28*16] = data_11_array[a19][b555][m555];
        end
    endgenerate
    generate 
        localparam integer b556 = 24;
        for (m556 = 0; m556 < 16; m556 = m556 + 1) 
        begin: inbit556
            assign data_11[m556 + b556*16 + a19*28*16] = data_11_array[a19][b556][m556];
        end
    endgenerate
    generate 
        localparam integer b557 = 25;
        for (m557 = 0; m557 < 16; m557 = m557 + 1) 
        begin: inbit557
            assign data_11[m557 + b557*16 + a19*28*16] = data_11_array[a19][b557][m557];
        end
    endgenerate
    generate 
        localparam integer b558 = 26;
        for (m558 = 0; m558 < 16; m558 = m558 + 1) 
        begin: inbit558
            assign data_11[m558 + b558*16 + a19*28*16] = data_11_array[a19][b558][m558];
        end
    endgenerate
    generate 
        localparam integer b559 = 27;
        for (m559 = 0; m559 < 16; m559 = m559 + 1) 
        begin: inbit559
            assign data_11[m559 + b559*16 + a19*28*16] = data_11_array[a19][b559][m559];
        end
    endgenerate
    localparam integer a20 = 20;
    generate 
        localparam integer b560 = 0;
        for (m560 = 0; m560 < 16; m560 = m560 + 1) 
        begin: inbit560
            assign data_11[m560 + b560*16 + a20*28*16] = data_11_array[a20][b560][m560];
        end
    endgenerate
    generate 
        localparam integer b561 = 1;
        for (m561 = 0; m561 < 16; m561 = m561 + 1) 
        begin: inbit561
            assign data_11[m561 + b561*16 + a20*28*16] = data_11_array[a20][b561][m561];
        end
    endgenerate
    generate 
        localparam integer b562 = 2;
        for (m562 = 0; m562 < 16; m562 = m562 + 1) 
        begin: inbit562
            assign data_11[m562 + b562*16 + a20*28*16] = data_11_array[a20][b562][m562];
        end
    endgenerate
    generate 
        localparam integer b563 = 3;
        for (m563 = 0; m563 < 16; m563 = m563 + 1) 
        begin: inbit563
            assign data_11[m563 + b563*16 + a20*28*16] = data_11_array[a20][b563][m563];
        end
    endgenerate
    generate 
        localparam integer b564 = 4;
        for (m564 = 0; m564 < 16; m564 = m564 + 1) 
        begin: inbit564
            assign data_11[m564 + b564*16 + a20*28*16] = data_11_array[a20][b564][m564];
        end
    endgenerate
    generate 
        localparam integer b565 = 5;
        for (m565 = 0; m565 < 16; m565 = m565 + 1) 
        begin: inbit565
            assign data_11[m565 + b565*16 + a20*28*16] = data_11_array[a20][b565][m565];
        end
    endgenerate
    generate 
        localparam integer b566 = 6;
        for (m566 = 0; m566 < 16; m566 = m566 + 1) 
        begin: inbit566
            assign data_11[m566 + b566*16 + a20*28*16] = data_11_array[a20][b566][m566];
        end
    endgenerate
    generate 
        localparam integer b567 = 7;
        for (m567 = 0; m567 < 16; m567 = m567 + 1) 
        begin: inbit567
            assign data_11[m567 + b567*16 + a20*28*16] = data_11_array[a20][b567][m567];
        end
    endgenerate
    generate 
        localparam integer b568 = 8;
        for (m568 = 0; m568 < 16; m568 = m568 + 1) 
        begin: inbit568
            assign data_11[m568 + b568*16 + a20*28*16] = data_11_array[a20][b568][m568];
        end
    endgenerate
    generate 
        localparam integer b569 = 9;
        for (m569 = 0; m569 < 16; m569 = m569 + 1) 
        begin: inbit569
            assign data_11[m569 + b569*16 + a20*28*16] = data_11_array[a20][b569][m569];
        end
    endgenerate
    generate 
        localparam integer b570 = 10;
        for (m570 = 0; m570 < 16; m570 = m570 + 1) 
        begin: inbit570
            assign data_11[m570 + b570*16 + a20*28*16] = data_11_array[a20][b570][m570];
        end
    endgenerate
    generate 
        localparam integer b571 = 11;
        for (m571 = 0; m571 < 16; m571 = m571 + 1) 
        begin: inbit571
            assign data_11[m571 + b571*16 + a20*28*16] = data_11_array[a20][b571][m571];
        end
    endgenerate
    generate 
        localparam integer b572 = 12;
        for (m572 = 0; m572 < 16; m572 = m572 + 1) 
        begin: inbit572
            assign data_11[m572 + b572*16 + a20*28*16] = data_11_array[a20][b572][m572];
        end
    endgenerate
    generate 
        localparam integer b573 = 13;
        for (m573 = 0; m573 < 16; m573 = m573 + 1) 
        begin: inbit573
            assign data_11[m573 + b573*16 + a20*28*16] = data_11_array[a20][b573][m573];
        end
    endgenerate
    generate 
        localparam integer b574 = 14;
        for (m574 = 0; m574 < 16; m574 = m574 + 1) 
        begin: inbit574
            assign data_11[m574 + b574*16 + a20*28*16] = data_11_array[a20][b574][m574];
        end
    endgenerate
    generate 
        localparam integer b575 = 15;
        for (m575 = 0; m575 < 16; m575 = m575 + 1) 
        begin: inbit575
            assign data_11[m575 + b575*16 + a20*28*16] = data_11_array[a20][b575][m575];
        end
    endgenerate
    generate 
        localparam integer b576 = 16;
        for (m576 = 0; m576 < 16; m576 = m576 + 1) 
        begin: inbit576
            assign data_11[m576 + b576*16 + a20*28*16] = data_11_array[a20][b576][m576];
        end
    endgenerate
    generate 
        localparam integer b577 = 17;
        for (m577 = 0; m577 < 16; m577 = m577 + 1) 
        begin: inbit577
            assign data_11[m577 + b577*16 + a20*28*16] = data_11_array[a20][b577][m577];
        end
    endgenerate
    generate 
        localparam integer b578 = 18;
        for (m578 = 0; m578 < 16; m578 = m578 + 1) 
        begin: inbit578
            assign data_11[m578 + b578*16 + a20*28*16] = data_11_array[a20][b578][m578];
        end
    endgenerate
    generate 
        localparam integer b579 = 19;
        for (m579 = 0; m579 < 16; m579 = m579 + 1) 
        begin: inbit579
            assign data_11[m579 + b579*16 + a20*28*16] = data_11_array[a20][b579][m579];
        end
    endgenerate
    generate 
        localparam integer b580 = 20;
        for (m580 = 0; m580 < 16; m580 = m580 + 1) 
        begin: inbit580
            assign data_11[m580 + b580*16 + a20*28*16] = data_11_array[a20][b580][m580];
        end
    endgenerate
    generate 
        localparam integer b581 = 21;
        for (m581 = 0; m581 < 16; m581 = m581 + 1) 
        begin: inbit581
            assign data_11[m581 + b581*16 + a20*28*16] = data_11_array[a20][b581][m581];
        end
    endgenerate
    generate 
        localparam integer b582 = 22;
        for (m582 = 0; m582 < 16; m582 = m582 + 1) 
        begin: inbit582
            assign data_11[m582 + b582*16 + a20*28*16] = data_11_array[a20][b582][m582];
        end
    endgenerate
    generate 
        localparam integer b583 = 23;
        for (m583 = 0; m583 < 16; m583 = m583 + 1) 
        begin: inbit583
            assign data_11[m583 + b583*16 + a20*28*16] = data_11_array[a20][b583][m583];
        end
    endgenerate
    generate 
        localparam integer b584 = 24;
        for (m584 = 0; m584 < 16; m584 = m584 + 1) 
        begin: inbit584
            assign data_11[m584 + b584*16 + a20*28*16] = data_11_array[a20][b584][m584];
        end
    endgenerate
    generate 
        localparam integer b585 = 25;
        for (m585 = 0; m585 < 16; m585 = m585 + 1) 
        begin: inbit585
            assign data_11[m585 + b585*16 + a20*28*16] = data_11_array[a20][b585][m585];
        end
    endgenerate
    generate 
        localparam integer b586 = 26;
        for (m586 = 0; m586 < 16; m586 = m586 + 1) 
        begin: inbit586
            assign data_11[m586 + b586*16 + a20*28*16] = data_11_array[a20][b586][m586];
        end
    endgenerate
    generate 
        localparam integer b587 = 27;
        for (m587 = 0; m587 < 16; m587 = m587 + 1) 
        begin: inbit587
            assign data_11[m587 + b587*16 + a20*28*16] = data_11_array[a20][b587][m587];
        end
    endgenerate
    localparam integer a21 = 21;
    generate 
        localparam integer b588 = 0;
        for (m588 = 0; m588 < 16; m588 = m588 + 1) 
        begin: inbit588
            assign data_11[m588 + b588*16 + a21*28*16] = data_11_array[a21][b588][m588];
        end
    endgenerate
    generate 
        localparam integer b589 = 1;
        for (m589 = 0; m589 < 16; m589 = m589 + 1) 
        begin: inbit589
            assign data_11[m589 + b589*16 + a21*28*16] = data_11_array[a21][b589][m589];
        end
    endgenerate
    generate 
        localparam integer b590 = 2;
        for (m590 = 0; m590 < 16; m590 = m590 + 1) 
        begin: inbit590
            assign data_11[m590 + b590*16 + a21*28*16] = data_11_array[a21][b590][m590];
        end
    endgenerate
    generate 
        localparam integer b591 = 3;
        for (m591 = 0; m591 < 16; m591 = m591 + 1) 
        begin: inbit591
            assign data_11[m591 + b591*16 + a21*28*16] = data_11_array[a21][b591][m591];
        end
    endgenerate
    generate 
        localparam integer b592 = 4;
        for (m592 = 0; m592 < 16; m592 = m592 + 1) 
        begin: inbit592
            assign data_11[m592 + b592*16 + a21*28*16] = data_11_array[a21][b592][m592];
        end
    endgenerate
    generate 
        localparam integer b593 = 5;
        for (m593 = 0; m593 < 16; m593 = m593 + 1) 
        begin: inbit593
            assign data_11[m593 + b593*16 + a21*28*16] = data_11_array[a21][b593][m593];
        end
    endgenerate
    generate 
        localparam integer b594 = 6;
        for (m594 = 0; m594 < 16; m594 = m594 + 1) 
        begin: inbit594
            assign data_11[m594 + b594*16 + a21*28*16] = data_11_array[a21][b594][m594];
        end
    endgenerate
    generate 
        localparam integer b595 = 7;
        for (m595 = 0; m595 < 16; m595 = m595 + 1) 
        begin: inbit595
            assign data_11[m595 + b595*16 + a21*28*16] = data_11_array[a21][b595][m595];
        end
    endgenerate
    generate 
        localparam integer b596 = 8;
        for (m596 = 0; m596 < 16; m596 = m596 + 1) 
        begin: inbit596
            assign data_11[m596 + b596*16 + a21*28*16] = data_11_array[a21][b596][m596];
        end
    endgenerate
    generate 
        localparam integer b597 = 9;
        for (m597 = 0; m597 < 16; m597 = m597 + 1) 
        begin: inbit597
            assign data_11[m597 + b597*16 + a21*28*16] = data_11_array[a21][b597][m597];
        end
    endgenerate
    generate 
        localparam integer b598 = 10;
        for (m598 = 0; m598 < 16; m598 = m598 + 1) 
        begin: inbit598
            assign data_11[m598 + b598*16 + a21*28*16] = data_11_array[a21][b598][m598];
        end
    endgenerate
    generate 
        localparam integer b599 = 11;
        for (m599 = 0; m599 < 16; m599 = m599 + 1) 
        begin: inbit599
            assign data_11[m599 + b599*16 + a21*28*16] = data_11_array[a21][b599][m599];
        end
    endgenerate
    generate 
        localparam integer b600 = 12;
        for (m600 = 0; m600 < 16; m600 = m600 + 1) 
        begin: inbit600
            assign data_11[m600 + b600*16 + a21*28*16] = data_11_array[a21][b600][m600];
        end
    endgenerate
    generate 
        localparam integer b601 = 13;
        for (m601 = 0; m601 < 16; m601 = m601 + 1) 
        begin: inbit601
            assign data_11[m601 + b601*16 + a21*28*16] = data_11_array[a21][b601][m601];
        end
    endgenerate
    generate 
        localparam integer b602 = 14;
        for (m602 = 0; m602 < 16; m602 = m602 + 1) 
        begin: inbit602
            assign data_11[m602 + b602*16 + a21*28*16] = data_11_array[a21][b602][m602];
        end
    endgenerate
    generate 
        localparam integer b603 = 15;
        for (m603 = 0; m603 < 16; m603 = m603 + 1) 
        begin: inbit603
            assign data_11[m603 + b603*16 + a21*28*16] = data_11_array[a21][b603][m603];
        end
    endgenerate
    generate 
        localparam integer b604 = 16;
        for (m604 = 0; m604 < 16; m604 = m604 + 1) 
        begin: inbit604
            assign data_11[m604 + b604*16 + a21*28*16] = data_11_array[a21][b604][m604];
        end
    endgenerate
    generate 
        localparam integer b605 = 17;
        for (m605 = 0; m605 < 16; m605 = m605 + 1) 
        begin: inbit605
            assign data_11[m605 + b605*16 + a21*28*16] = data_11_array[a21][b605][m605];
        end
    endgenerate
    generate 
        localparam integer b606 = 18;
        for (m606 = 0; m606 < 16; m606 = m606 + 1) 
        begin: inbit606
            assign data_11[m606 + b606*16 + a21*28*16] = data_11_array[a21][b606][m606];
        end
    endgenerate
    generate 
        localparam integer b607 = 19;
        for (m607 = 0; m607 < 16; m607 = m607 + 1) 
        begin: inbit607
            assign data_11[m607 + b607*16 + a21*28*16] = data_11_array[a21][b607][m607];
        end
    endgenerate
    generate 
        localparam integer b608 = 20;
        for (m608 = 0; m608 < 16; m608 = m608 + 1) 
        begin: inbit608
            assign data_11[m608 + b608*16 + a21*28*16] = data_11_array[a21][b608][m608];
        end
    endgenerate
    generate 
        localparam integer b609 = 21;
        for (m609 = 0; m609 < 16; m609 = m609 + 1) 
        begin: inbit609
            assign data_11[m609 + b609*16 + a21*28*16] = data_11_array[a21][b609][m609];
        end
    endgenerate
    generate 
        localparam integer b610 = 22;
        for (m610 = 0; m610 < 16; m610 = m610 + 1) 
        begin: inbit610
            assign data_11[m610 + b610*16 + a21*28*16] = data_11_array[a21][b610][m610];
        end
    endgenerate
    generate 
        localparam integer b611 = 23;
        for (m611 = 0; m611 < 16; m611 = m611 + 1) 
        begin: inbit611
            assign data_11[m611 + b611*16 + a21*28*16] = data_11_array[a21][b611][m611];
        end
    endgenerate
    generate 
        localparam integer b612 = 24;
        for (m612 = 0; m612 < 16; m612 = m612 + 1) 
        begin: inbit612
            assign data_11[m612 + b612*16 + a21*28*16] = data_11_array[a21][b612][m612];
        end
    endgenerate
    generate 
        localparam integer b613 = 25;
        for (m613 = 0; m613 < 16; m613 = m613 + 1) 
        begin: inbit613
            assign data_11[m613 + b613*16 + a21*28*16] = data_11_array[a21][b613][m613];
        end
    endgenerate
    generate 
        localparam integer b614 = 26;
        for (m614 = 0; m614 < 16; m614 = m614 + 1) 
        begin: inbit614
            assign data_11[m614 + b614*16 + a21*28*16] = data_11_array[a21][b614][m614];
        end
    endgenerate
    generate 
        localparam integer b615 = 27;
        for (m615 = 0; m615 < 16; m615 = m615 + 1) 
        begin: inbit615
            assign data_11[m615 + b615*16 + a21*28*16] = data_11_array[a21][b615][m615];
        end
    endgenerate
    localparam integer a22 = 22;
    generate 
        localparam integer b616 = 0;
        for (m616 = 0; m616 < 16; m616 = m616 + 1) 
        begin: inbit616
            assign data_11[m616 + b616*16 + a22*28*16] = data_11_array[a22][b616][m616];
        end
    endgenerate
    generate 
        localparam integer b617 = 1;
        for (m617 = 0; m617 < 16; m617 = m617 + 1) 
        begin: inbit617
            assign data_11[m617 + b617*16 + a22*28*16] = data_11_array[a22][b617][m617];
        end
    endgenerate
    generate 
        localparam integer b618 = 2;
        for (m618 = 0; m618 < 16; m618 = m618 + 1) 
        begin: inbit618
            assign data_11[m618 + b618*16 + a22*28*16] = data_11_array[a22][b618][m618];
        end
    endgenerate
    generate 
        localparam integer b619 = 3;
        for (m619 = 0; m619 < 16; m619 = m619 + 1) 
        begin: inbit619
            assign data_11[m619 + b619*16 + a22*28*16] = data_11_array[a22][b619][m619];
        end
    endgenerate
    generate 
        localparam integer b620 = 4;
        for (m620 = 0; m620 < 16; m620 = m620 + 1) 
        begin: inbit620
            assign data_11[m620 + b620*16 + a22*28*16] = data_11_array[a22][b620][m620];
        end
    endgenerate
    generate 
        localparam integer b621 = 5;
        for (m621 = 0; m621 < 16; m621 = m621 + 1) 
        begin: inbit621
            assign data_11[m621 + b621*16 + a22*28*16] = data_11_array[a22][b621][m621];
        end
    endgenerate
    generate 
        localparam integer b622 = 6;
        for (m622 = 0; m622 < 16; m622 = m622 + 1) 
        begin: inbit622
            assign data_11[m622 + b622*16 + a22*28*16] = data_11_array[a22][b622][m622];
        end
    endgenerate
    generate 
        localparam integer b623 = 7;
        for (m623 = 0; m623 < 16; m623 = m623 + 1) 
        begin: inbit623
            assign data_11[m623 + b623*16 + a22*28*16] = data_11_array[a22][b623][m623];
        end
    endgenerate
    generate 
        localparam integer b624 = 8;
        for (m624 = 0; m624 < 16; m624 = m624 + 1) 
        begin: inbit624
            assign data_11[m624 + b624*16 + a22*28*16] = data_11_array[a22][b624][m624];
        end
    endgenerate
    generate 
        localparam integer b625 = 9;
        for (m625 = 0; m625 < 16; m625 = m625 + 1) 
        begin: inbit625
            assign data_11[m625 + b625*16 + a22*28*16] = data_11_array[a22][b625][m625];
        end
    endgenerate
    generate 
        localparam integer b626 = 10;
        for (m626 = 0; m626 < 16; m626 = m626 + 1) 
        begin: inbit626
            assign data_11[m626 + b626*16 + a22*28*16] = data_11_array[a22][b626][m626];
        end
    endgenerate
    generate 
        localparam integer b627 = 11;
        for (m627 = 0; m627 < 16; m627 = m627 + 1) 
        begin: inbit627
            assign data_11[m627 + b627*16 + a22*28*16] = data_11_array[a22][b627][m627];
        end
    endgenerate
    generate 
        localparam integer b628 = 12;
        for (m628 = 0; m628 < 16; m628 = m628 + 1) 
        begin: inbit628
            assign data_11[m628 + b628*16 + a22*28*16] = data_11_array[a22][b628][m628];
        end
    endgenerate
    generate 
        localparam integer b629 = 13;
        for (m629 = 0; m629 < 16; m629 = m629 + 1) 
        begin: inbit629
            assign data_11[m629 + b629*16 + a22*28*16] = data_11_array[a22][b629][m629];
        end
    endgenerate
    generate 
        localparam integer b630 = 14;
        for (m630 = 0; m630 < 16; m630 = m630 + 1) 
        begin: inbit630
            assign data_11[m630 + b630*16 + a22*28*16] = data_11_array[a22][b630][m630];
        end
    endgenerate
    generate 
        localparam integer b631 = 15;
        for (m631 = 0; m631 < 16; m631 = m631 + 1) 
        begin: inbit631
            assign data_11[m631 + b631*16 + a22*28*16] = data_11_array[a22][b631][m631];
        end
    endgenerate
    generate 
        localparam integer b632 = 16;
        for (m632 = 0; m632 < 16; m632 = m632 + 1) 
        begin: inbit632
            assign data_11[m632 + b632*16 + a22*28*16] = data_11_array[a22][b632][m632];
        end
    endgenerate
    generate 
        localparam integer b633 = 17;
        for (m633 = 0; m633 < 16; m633 = m633 + 1) 
        begin: inbit633
            assign data_11[m633 + b633*16 + a22*28*16] = data_11_array[a22][b633][m633];
        end
    endgenerate
    generate 
        localparam integer b634 = 18;
        for (m634 = 0; m634 < 16; m634 = m634 + 1) 
        begin: inbit634
            assign data_11[m634 + b634*16 + a22*28*16] = data_11_array[a22][b634][m634];
        end
    endgenerate
    generate 
        localparam integer b635 = 19;
        for (m635 = 0; m635 < 16; m635 = m635 + 1) 
        begin: inbit635
            assign data_11[m635 + b635*16 + a22*28*16] = data_11_array[a22][b635][m635];
        end
    endgenerate
    generate 
        localparam integer b636 = 20;
        for (m636 = 0; m636 < 16; m636 = m636 + 1) 
        begin: inbit636
            assign data_11[m636 + b636*16 + a22*28*16] = data_11_array[a22][b636][m636];
        end
    endgenerate
    generate 
        localparam integer b637 = 21;
        for (m637 = 0; m637 < 16; m637 = m637 + 1) 
        begin: inbit637
            assign data_11[m637 + b637*16 + a22*28*16] = data_11_array[a22][b637][m637];
        end
    endgenerate
    generate 
        localparam integer b638 = 22;
        for (m638 = 0; m638 < 16; m638 = m638 + 1) 
        begin: inbit638
            assign data_11[m638 + b638*16 + a22*28*16] = data_11_array[a22][b638][m638];
        end
    endgenerate
    generate 
        localparam integer b639 = 23;
        for (m639 = 0; m639 < 16; m639 = m639 + 1) 
        begin: inbit639
            assign data_11[m639 + b639*16 + a22*28*16] = data_11_array[a22][b639][m639];
        end
    endgenerate
    generate 
        localparam integer b640 = 24;
        for (m640 = 0; m640 < 16; m640 = m640 + 1) 
        begin: inbit640
            assign data_11[m640 + b640*16 + a22*28*16] = data_11_array[a22][b640][m640];
        end
    endgenerate
    generate 
        localparam integer b641 = 25;
        for (m641 = 0; m641 < 16; m641 = m641 + 1) 
        begin: inbit641
            assign data_11[m641 + b641*16 + a22*28*16] = data_11_array[a22][b641][m641];
        end
    endgenerate
    generate 
        localparam integer b642 = 26;
        for (m642 = 0; m642 < 16; m642 = m642 + 1) 
        begin: inbit642
            assign data_11[m642 + b642*16 + a22*28*16] = data_11_array[a22][b642][m642];
        end
    endgenerate
    generate 
        localparam integer b643 = 27;
        for (m643 = 0; m643 < 16; m643 = m643 + 1) 
        begin: inbit643
            assign data_11[m643 + b643*16 + a22*28*16] = data_11_array[a22][b643][m643];
        end
    endgenerate
    localparam integer a23 = 23;
    generate 
        localparam integer b644 = 0;
        for (m644 = 0; m644 < 16; m644 = m644 + 1) 
        begin: inbit644
            assign data_11[m644 + b644*16 + a23*28*16] = data_11_array[a23][b644][m644];
        end
    endgenerate
    generate 
        localparam integer b645 = 1;
        for (m645 = 0; m645 < 16; m645 = m645 + 1) 
        begin: inbit645
            assign data_11[m645 + b645*16 + a23*28*16] = data_11_array[a23][b645][m645];
        end
    endgenerate
    generate 
        localparam integer b646 = 2;
        for (m646 = 0; m646 < 16; m646 = m646 + 1) 
        begin: inbit646
            assign data_11[m646 + b646*16 + a23*28*16] = data_11_array[a23][b646][m646];
        end
    endgenerate
    generate 
        localparam integer b647 = 3;
        for (m647 = 0; m647 < 16; m647 = m647 + 1) 
        begin: inbit647
            assign data_11[m647 + b647*16 + a23*28*16] = data_11_array[a23][b647][m647];
        end
    endgenerate
    generate 
        localparam integer b648 = 4;
        for (m648 = 0; m648 < 16; m648 = m648 + 1) 
        begin: inbit648
            assign data_11[m648 + b648*16 + a23*28*16] = data_11_array[a23][b648][m648];
        end
    endgenerate
    generate 
        localparam integer b649 = 5;
        for (m649 = 0; m649 < 16; m649 = m649 + 1) 
        begin: inbit649
            assign data_11[m649 + b649*16 + a23*28*16] = data_11_array[a23][b649][m649];
        end
    endgenerate
    generate 
        localparam integer b650 = 6;
        for (m650 = 0; m650 < 16; m650 = m650 + 1) 
        begin: inbit650
            assign data_11[m650 + b650*16 + a23*28*16] = data_11_array[a23][b650][m650];
        end
    endgenerate
    generate 
        localparam integer b651 = 7;
        for (m651 = 0; m651 < 16; m651 = m651 + 1) 
        begin: inbit651
            assign data_11[m651 + b651*16 + a23*28*16] = data_11_array[a23][b651][m651];
        end
    endgenerate
    generate 
        localparam integer b652 = 8;
        for (m652 = 0; m652 < 16; m652 = m652 + 1) 
        begin: inbit652
            assign data_11[m652 + b652*16 + a23*28*16] = data_11_array[a23][b652][m652];
        end
    endgenerate
    generate 
        localparam integer b653 = 9;
        for (m653 = 0; m653 < 16; m653 = m653 + 1) 
        begin: inbit653
            assign data_11[m653 + b653*16 + a23*28*16] = data_11_array[a23][b653][m653];
        end
    endgenerate
    generate 
        localparam integer b654 = 10;
        for (m654 = 0; m654 < 16; m654 = m654 + 1) 
        begin: inbit654
            assign data_11[m654 + b654*16 + a23*28*16] = data_11_array[a23][b654][m654];
        end
    endgenerate
    generate 
        localparam integer b655 = 11;
        for (m655 = 0; m655 < 16; m655 = m655 + 1) 
        begin: inbit655
            assign data_11[m655 + b655*16 + a23*28*16] = data_11_array[a23][b655][m655];
        end
    endgenerate
    generate 
        localparam integer b656 = 12;
        for (m656 = 0; m656 < 16; m656 = m656 + 1) 
        begin: inbit656
            assign data_11[m656 + b656*16 + a23*28*16] = data_11_array[a23][b656][m656];
        end
    endgenerate
    generate 
        localparam integer b657 = 13;
        for (m657 = 0; m657 < 16; m657 = m657 + 1) 
        begin: inbit657
            assign data_11[m657 + b657*16 + a23*28*16] = data_11_array[a23][b657][m657];
        end
    endgenerate
    generate 
        localparam integer b658 = 14;
        for (m658 = 0; m658 < 16; m658 = m658 + 1) 
        begin: inbit658
            assign data_11[m658 + b658*16 + a23*28*16] = data_11_array[a23][b658][m658];
        end
    endgenerate
    generate 
        localparam integer b659 = 15;
        for (m659 = 0; m659 < 16; m659 = m659 + 1) 
        begin: inbit659
            assign data_11[m659 + b659*16 + a23*28*16] = data_11_array[a23][b659][m659];
        end
    endgenerate
    generate 
        localparam integer b660 = 16;
        for (m660 = 0; m660 < 16; m660 = m660 + 1) 
        begin: inbit660
            assign data_11[m660 + b660*16 + a23*28*16] = data_11_array[a23][b660][m660];
        end
    endgenerate
    generate 
        localparam integer b661 = 17;
        for (m661 = 0; m661 < 16; m661 = m661 + 1) 
        begin: inbit661
            assign data_11[m661 + b661*16 + a23*28*16] = data_11_array[a23][b661][m661];
        end
    endgenerate
    generate 
        localparam integer b662 = 18;
        for (m662 = 0; m662 < 16; m662 = m662 + 1) 
        begin: inbit662
            assign data_11[m662 + b662*16 + a23*28*16] = data_11_array[a23][b662][m662];
        end
    endgenerate
    generate 
        localparam integer b663 = 19;
        for (m663 = 0; m663 < 16; m663 = m663 + 1) 
        begin: inbit663
            assign data_11[m663 + b663*16 + a23*28*16] = data_11_array[a23][b663][m663];
        end
    endgenerate
    generate 
        localparam integer b664 = 20;
        for (m664 = 0; m664 < 16; m664 = m664 + 1) 
        begin: inbit664
            assign data_11[m664 + b664*16 + a23*28*16] = data_11_array[a23][b664][m664];
        end
    endgenerate
    generate 
        localparam integer b665 = 21;
        for (m665 = 0; m665 < 16; m665 = m665 + 1) 
        begin: inbit665
            assign data_11[m665 + b665*16 + a23*28*16] = data_11_array[a23][b665][m665];
        end
    endgenerate
    generate 
        localparam integer b666 = 22;
        for (m666 = 0; m666 < 16; m666 = m666 + 1) 
        begin: inbit666
            assign data_11[m666 + b666*16 + a23*28*16] = data_11_array[a23][b666][m666];
        end
    endgenerate
    generate 
        localparam integer b667 = 23;
        for (m667 = 0; m667 < 16; m667 = m667 + 1) 
        begin: inbit667
            assign data_11[m667 + b667*16 + a23*28*16] = data_11_array[a23][b667][m667];
        end
    endgenerate
    generate 
        localparam integer b668 = 24;
        for (m668 = 0; m668 < 16; m668 = m668 + 1) 
        begin: inbit668
            assign data_11[m668 + b668*16 + a23*28*16] = data_11_array[a23][b668][m668];
        end
    endgenerate
    generate 
        localparam integer b669 = 25;
        for (m669 = 0; m669 < 16; m669 = m669 + 1) 
        begin: inbit669
            assign data_11[m669 + b669*16 + a23*28*16] = data_11_array[a23][b669][m669];
        end
    endgenerate
    generate 
        localparam integer b670 = 26;
        for (m670 = 0; m670 < 16; m670 = m670 + 1) 
        begin: inbit670
            assign data_11[m670 + b670*16 + a23*28*16] = data_11_array[a23][b670][m670];
        end
    endgenerate
    generate 
        localparam integer b671 = 27;
        for (m671 = 0; m671 < 16; m671 = m671 + 1) 
        begin: inbit671
            assign data_11[m671 + b671*16 + a23*28*16] = data_11_array[a23][b671][m671];
        end
    endgenerate
    localparam integer a24 = 24;
    generate 
        localparam integer b672 = 0;
        for (m672 = 0; m672 < 16; m672 = m672 + 1) 
        begin: inbit672
            assign data_11[m672 + b672*16 + a24*28*16] = data_11_array[a24][b672][m672];
        end
    endgenerate
    generate 
        localparam integer b673 = 1;
        for (m673 = 0; m673 < 16; m673 = m673 + 1) 
        begin: inbit673
            assign data_11[m673 + b673*16 + a24*28*16] = data_11_array[a24][b673][m673];
        end
    endgenerate
    generate 
        localparam integer b674 = 2;
        for (m674 = 0; m674 < 16; m674 = m674 + 1) 
        begin: inbit674
            assign data_11[m674 + b674*16 + a24*28*16] = data_11_array[a24][b674][m674];
        end
    endgenerate
    generate 
        localparam integer b675 = 3;
        for (m675 = 0; m675 < 16; m675 = m675 + 1) 
        begin: inbit675
            assign data_11[m675 + b675*16 + a24*28*16] = data_11_array[a24][b675][m675];
        end
    endgenerate
    generate 
        localparam integer b676 = 4;
        for (m676 = 0; m676 < 16; m676 = m676 + 1) 
        begin: inbit676
            assign data_11[m676 + b676*16 + a24*28*16] = data_11_array[a24][b676][m676];
        end
    endgenerate
    generate 
        localparam integer b677 = 5;
        for (m677 = 0; m677 < 16; m677 = m677 + 1) 
        begin: inbit677
            assign data_11[m677 + b677*16 + a24*28*16] = data_11_array[a24][b677][m677];
        end
    endgenerate
    generate 
        localparam integer b678 = 6;
        for (m678 = 0; m678 < 16; m678 = m678 + 1) 
        begin: inbit678
            assign data_11[m678 + b678*16 + a24*28*16] = data_11_array[a24][b678][m678];
        end
    endgenerate
    generate 
        localparam integer b679 = 7;
        for (m679 = 0; m679 < 16; m679 = m679 + 1) 
        begin: inbit679
            assign data_11[m679 + b679*16 + a24*28*16] = data_11_array[a24][b679][m679];
        end
    endgenerate
    generate 
        localparam integer b680 = 8;
        for (m680 = 0; m680 < 16; m680 = m680 + 1) 
        begin: inbit680
            assign data_11[m680 + b680*16 + a24*28*16] = data_11_array[a24][b680][m680];
        end
    endgenerate
    generate 
        localparam integer b681 = 9;
        for (m681 = 0; m681 < 16; m681 = m681 + 1) 
        begin: inbit681
            assign data_11[m681 + b681*16 + a24*28*16] = data_11_array[a24][b681][m681];
        end
    endgenerate
    generate 
        localparam integer b682 = 10;
        for (m682 = 0; m682 < 16; m682 = m682 + 1) 
        begin: inbit682
            assign data_11[m682 + b682*16 + a24*28*16] = data_11_array[a24][b682][m682];
        end
    endgenerate
    generate 
        localparam integer b683 = 11;
        for (m683 = 0; m683 < 16; m683 = m683 + 1) 
        begin: inbit683
            assign data_11[m683 + b683*16 + a24*28*16] = data_11_array[a24][b683][m683];
        end
    endgenerate
    generate 
        localparam integer b684 = 12;
        for (m684 = 0; m684 < 16; m684 = m684 + 1) 
        begin: inbit684
            assign data_11[m684 + b684*16 + a24*28*16] = data_11_array[a24][b684][m684];
        end
    endgenerate
    generate 
        localparam integer b685 = 13;
        for (m685 = 0; m685 < 16; m685 = m685 + 1) 
        begin: inbit685
            assign data_11[m685 + b685*16 + a24*28*16] = data_11_array[a24][b685][m685];
        end
    endgenerate
    generate 
        localparam integer b686 = 14;
        for (m686 = 0; m686 < 16; m686 = m686 + 1) 
        begin: inbit686
            assign data_11[m686 + b686*16 + a24*28*16] = data_11_array[a24][b686][m686];
        end
    endgenerate
    generate 
        localparam integer b687 = 15;
        for (m687 = 0; m687 < 16; m687 = m687 + 1) 
        begin: inbit687
            assign data_11[m687 + b687*16 + a24*28*16] = data_11_array[a24][b687][m687];
        end
    endgenerate
    generate 
        localparam integer b688 = 16;
        for (m688 = 0; m688 < 16; m688 = m688 + 1) 
        begin: inbit688
            assign data_11[m688 + b688*16 + a24*28*16] = data_11_array[a24][b688][m688];
        end
    endgenerate
    generate 
        localparam integer b689 = 17;
        for (m689 = 0; m689 < 16; m689 = m689 + 1) 
        begin: inbit689
            assign data_11[m689 + b689*16 + a24*28*16] = data_11_array[a24][b689][m689];
        end
    endgenerate
    generate 
        localparam integer b690 = 18;
        for (m690 = 0; m690 < 16; m690 = m690 + 1) 
        begin: inbit690
            assign data_11[m690 + b690*16 + a24*28*16] = data_11_array[a24][b690][m690];
        end
    endgenerate
    generate 
        localparam integer b691 = 19;
        for (m691 = 0; m691 < 16; m691 = m691 + 1) 
        begin: inbit691
            assign data_11[m691 + b691*16 + a24*28*16] = data_11_array[a24][b691][m691];
        end
    endgenerate
    generate 
        localparam integer b692 = 20;
        for (m692 = 0; m692 < 16; m692 = m692 + 1) 
        begin: inbit692
            assign data_11[m692 + b692*16 + a24*28*16] = data_11_array[a24][b692][m692];
        end
    endgenerate
    generate 
        localparam integer b693 = 21;
        for (m693 = 0; m693 < 16; m693 = m693 + 1) 
        begin: inbit693
            assign data_11[m693 + b693*16 + a24*28*16] = data_11_array[a24][b693][m693];
        end
    endgenerate
    generate 
        localparam integer b694 = 22;
        for (m694 = 0; m694 < 16; m694 = m694 + 1) 
        begin: inbit694
            assign data_11[m694 + b694*16 + a24*28*16] = data_11_array[a24][b694][m694];
        end
    endgenerate
    generate 
        localparam integer b695 = 23;
        for (m695 = 0; m695 < 16; m695 = m695 + 1) 
        begin: inbit695
            assign data_11[m695 + b695*16 + a24*28*16] = data_11_array[a24][b695][m695];
        end
    endgenerate
    generate 
        localparam integer b696 = 24;
        for (m696 = 0; m696 < 16; m696 = m696 + 1) 
        begin: inbit696
            assign data_11[m696 + b696*16 + a24*28*16] = data_11_array[a24][b696][m696];
        end
    endgenerate
    generate 
        localparam integer b697 = 25;
        for (m697 = 0; m697 < 16; m697 = m697 + 1) 
        begin: inbit697
            assign data_11[m697 + b697*16 + a24*28*16] = data_11_array[a24][b697][m697];
        end
    endgenerate
    generate 
        localparam integer b698 = 26;
        for (m698 = 0; m698 < 16; m698 = m698 + 1) 
        begin: inbit698
            assign data_11[m698 + b698*16 + a24*28*16] = data_11_array[a24][b698][m698];
        end
    endgenerate
    generate 
        localparam integer b699 = 27;
        for (m699 = 0; m699 < 16; m699 = m699 + 1) 
        begin: inbit699
            assign data_11[m699 + b699*16 + a24*28*16] = data_11_array[a24][b699][m699];
        end
    endgenerate
    localparam integer a25 = 25;
    generate 
        localparam integer b700 = 0;
        for (m700 = 0; m700 < 16; m700 = m700 + 1) 
        begin: inbit700
            assign data_11[m700 + b700*16 + a25*28*16] = data_11_array[a25][b700][m700];
        end
    endgenerate
    generate 
        localparam integer b701 = 1;
        for (m701 = 0; m701 < 16; m701 = m701 + 1) 
        begin: inbit701
            assign data_11[m701 + b701*16 + a25*28*16] = data_11_array[a25][b701][m701];
        end
    endgenerate
    generate 
        localparam integer b702 = 2;
        for (m702 = 0; m702 < 16; m702 = m702 + 1) 
        begin: inbit702
            assign data_11[m702 + b702*16 + a25*28*16] = data_11_array[a25][b702][m702];
        end
    endgenerate
    generate 
        localparam integer b703 = 3;
        for (m703 = 0; m703 < 16; m703 = m703 + 1) 
        begin: inbit703
            assign data_11[m703 + b703*16 + a25*28*16] = data_11_array[a25][b703][m703];
        end
    endgenerate
    generate 
        localparam integer b704 = 4;
        for (m704 = 0; m704 < 16; m704 = m704 + 1) 
        begin: inbit704
            assign data_11[m704 + b704*16 + a25*28*16] = data_11_array[a25][b704][m704];
        end
    endgenerate
    generate 
        localparam integer b705 = 5;
        for (m705 = 0; m705 < 16; m705 = m705 + 1) 
        begin: inbit705
            assign data_11[m705 + b705*16 + a25*28*16] = data_11_array[a25][b705][m705];
        end
    endgenerate
    generate 
        localparam integer b706 = 6;
        for (m706 = 0; m706 < 16; m706 = m706 + 1) 
        begin: inbit706
            assign data_11[m706 + b706*16 + a25*28*16] = data_11_array[a25][b706][m706];
        end
    endgenerate
    generate 
        localparam integer b707 = 7;
        for (m707 = 0; m707 < 16; m707 = m707 + 1) 
        begin: inbit707
            assign data_11[m707 + b707*16 + a25*28*16] = data_11_array[a25][b707][m707];
        end
    endgenerate
    generate 
        localparam integer b708 = 8;
        for (m708 = 0; m708 < 16; m708 = m708 + 1) 
        begin: inbit708
            assign data_11[m708 + b708*16 + a25*28*16] = data_11_array[a25][b708][m708];
        end
    endgenerate
    generate 
        localparam integer b709 = 9;
        for (m709 = 0; m709 < 16; m709 = m709 + 1) 
        begin: inbit709
            assign data_11[m709 + b709*16 + a25*28*16] = data_11_array[a25][b709][m709];
        end
    endgenerate
    generate 
        localparam integer b710 = 10;
        for (m710 = 0; m710 < 16; m710 = m710 + 1) 
        begin: inbit710
            assign data_11[m710 + b710*16 + a25*28*16] = data_11_array[a25][b710][m710];
        end
    endgenerate
    generate 
        localparam integer b711 = 11;
        for (m711 = 0; m711 < 16; m711 = m711 + 1) 
        begin: inbit711
            assign data_11[m711 + b711*16 + a25*28*16] = data_11_array[a25][b711][m711];
        end
    endgenerate
    generate 
        localparam integer b712 = 12;
        for (m712 = 0; m712 < 16; m712 = m712 + 1) 
        begin: inbit712
            assign data_11[m712 + b712*16 + a25*28*16] = data_11_array[a25][b712][m712];
        end
    endgenerate
    generate 
        localparam integer b713 = 13;
        for (m713 = 0; m713 < 16; m713 = m713 + 1) 
        begin: inbit713
            assign data_11[m713 + b713*16 + a25*28*16] = data_11_array[a25][b713][m713];
        end
    endgenerate
    generate 
        localparam integer b714 = 14;
        for (m714 = 0; m714 < 16; m714 = m714 + 1) 
        begin: inbit714
            assign data_11[m714 + b714*16 + a25*28*16] = data_11_array[a25][b714][m714];
        end
    endgenerate
    generate 
        localparam integer b715 = 15;
        for (m715 = 0; m715 < 16; m715 = m715 + 1) 
        begin: inbit715
            assign data_11[m715 + b715*16 + a25*28*16] = data_11_array[a25][b715][m715];
        end
    endgenerate
    generate 
        localparam integer b716 = 16;
        for (m716 = 0; m716 < 16; m716 = m716 + 1) 
        begin: inbit716
            assign data_11[m716 + b716*16 + a25*28*16] = data_11_array[a25][b716][m716];
        end
    endgenerate
    generate 
        localparam integer b717 = 17;
        for (m717 = 0; m717 < 16; m717 = m717 + 1) 
        begin: inbit717
            assign data_11[m717 + b717*16 + a25*28*16] = data_11_array[a25][b717][m717];
        end
    endgenerate
    generate 
        localparam integer b718 = 18;
        for (m718 = 0; m718 < 16; m718 = m718 + 1) 
        begin: inbit718
            assign data_11[m718 + b718*16 + a25*28*16] = data_11_array[a25][b718][m718];
        end
    endgenerate
    generate 
        localparam integer b719 = 19;
        for (m719 = 0; m719 < 16; m719 = m719 + 1) 
        begin: inbit719
            assign data_11[m719 + b719*16 + a25*28*16] = data_11_array[a25][b719][m719];
        end
    endgenerate
    generate 
        localparam integer b720 = 20;
        for (m720 = 0; m720 < 16; m720 = m720 + 1) 
        begin: inbit720
            assign data_11[m720 + b720*16 + a25*28*16] = data_11_array[a25][b720][m720];
        end
    endgenerate
    generate 
        localparam integer b721 = 21;
        for (m721 = 0; m721 < 16; m721 = m721 + 1) 
        begin: inbit721
            assign data_11[m721 + b721*16 + a25*28*16] = data_11_array[a25][b721][m721];
        end
    endgenerate
    generate 
        localparam integer b722 = 22;
        for (m722 = 0; m722 < 16; m722 = m722 + 1) 
        begin: inbit722
            assign data_11[m722 + b722*16 + a25*28*16] = data_11_array[a25][b722][m722];
        end
    endgenerate
    generate 
        localparam integer b723 = 23;
        for (m723 = 0; m723 < 16; m723 = m723 + 1) 
        begin: inbit723
            assign data_11[m723 + b723*16 + a25*28*16] = data_11_array[a25][b723][m723];
        end
    endgenerate
    generate 
        localparam integer b724 = 24;
        for (m724 = 0; m724 < 16; m724 = m724 + 1) 
        begin: inbit724
            assign data_11[m724 + b724*16 + a25*28*16] = data_11_array[a25][b724][m724];
        end
    endgenerate
    generate 
        localparam integer b725 = 25;
        for (m725 = 0; m725 < 16; m725 = m725 + 1) 
        begin: inbit725
            assign data_11[m725 + b725*16 + a25*28*16] = data_11_array[a25][b725][m725];
        end
    endgenerate
    generate 
        localparam integer b726 = 26;
        for (m726 = 0; m726 < 16; m726 = m726 + 1) 
        begin: inbit726
            assign data_11[m726 + b726*16 + a25*28*16] = data_11_array[a25][b726][m726];
        end
    endgenerate
    generate 
        localparam integer b727 = 27;
        for (m727 = 0; m727 < 16; m727 = m727 + 1) 
        begin: inbit727
            assign data_11[m727 + b727*16 + a25*28*16] = data_11_array[a25][b727][m727];
        end
    endgenerate
    localparam integer a26 = 26;
    generate 
        localparam integer b728 = 0;
        for (m728 = 0; m728 < 16; m728 = m728 + 1) 
        begin: inbit728
            assign data_11[m728 + b728*16 + a26*28*16] = data_11_array[a26][b728][m728];
        end
    endgenerate
    generate 
        localparam integer b729 = 1;
        for (m729 = 0; m729 < 16; m729 = m729 + 1) 
        begin: inbit729
            assign data_11[m729 + b729*16 + a26*28*16] = data_11_array[a26][b729][m729];
        end
    endgenerate
    generate 
        localparam integer b730 = 2;
        for (m730 = 0; m730 < 16; m730 = m730 + 1) 
        begin: inbit730
            assign data_11[m730 + b730*16 + a26*28*16] = data_11_array[a26][b730][m730];
        end
    endgenerate
    generate 
        localparam integer b731 = 3;
        for (m731 = 0; m731 < 16; m731 = m731 + 1) 
        begin: inbit731
            assign data_11[m731 + b731*16 + a26*28*16] = data_11_array[a26][b731][m731];
        end
    endgenerate
    generate 
        localparam integer b732 = 4;
        for (m732 = 0; m732 < 16; m732 = m732 + 1) 
        begin: inbit732
            assign data_11[m732 + b732*16 + a26*28*16] = data_11_array[a26][b732][m732];
        end
    endgenerate
    generate 
        localparam integer b733 = 5;
        for (m733 = 0; m733 < 16; m733 = m733 + 1) 
        begin: inbit733
            assign data_11[m733 + b733*16 + a26*28*16] = data_11_array[a26][b733][m733];
        end
    endgenerate
    generate 
        localparam integer b734 = 6;
        for (m734 = 0; m734 < 16; m734 = m734 + 1) 
        begin: inbit734
            assign data_11[m734 + b734*16 + a26*28*16] = data_11_array[a26][b734][m734];
        end
    endgenerate
    generate 
        localparam integer b735 = 7;
        for (m735 = 0; m735 < 16; m735 = m735 + 1) 
        begin: inbit735
            assign data_11[m735 + b735*16 + a26*28*16] = data_11_array[a26][b735][m735];
        end
    endgenerate
    generate 
        localparam integer b736 = 8;
        for (m736 = 0; m736 < 16; m736 = m736 + 1) 
        begin: inbit736
            assign data_11[m736 + b736*16 + a26*28*16] = data_11_array[a26][b736][m736];
        end
    endgenerate
    generate 
        localparam integer b737 = 9;
        for (m737 = 0; m737 < 16; m737 = m737 + 1) 
        begin: inbit737
            assign data_11[m737 + b737*16 + a26*28*16] = data_11_array[a26][b737][m737];
        end
    endgenerate
    generate 
        localparam integer b738 = 10;
        for (m738 = 0; m738 < 16; m738 = m738 + 1) 
        begin: inbit738
            assign data_11[m738 + b738*16 + a26*28*16] = data_11_array[a26][b738][m738];
        end
    endgenerate
    generate 
        localparam integer b739 = 11;
        for (m739 = 0; m739 < 16; m739 = m739 + 1) 
        begin: inbit739
            assign data_11[m739 + b739*16 + a26*28*16] = data_11_array[a26][b739][m739];
        end
    endgenerate
    generate 
        localparam integer b740 = 12;
        for (m740 = 0; m740 < 16; m740 = m740 + 1) 
        begin: inbit740
            assign data_11[m740 + b740*16 + a26*28*16] = data_11_array[a26][b740][m740];
        end
    endgenerate
    generate 
        localparam integer b741 = 13;
        for (m741 = 0; m741 < 16; m741 = m741 + 1) 
        begin: inbit741
            assign data_11[m741 + b741*16 + a26*28*16] = data_11_array[a26][b741][m741];
        end
    endgenerate
    generate 
        localparam integer b742 = 14;
        for (m742 = 0; m742 < 16; m742 = m742 + 1) 
        begin: inbit742
            assign data_11[m742 + b742*16 + a26*28*16] = data_11_array[a26][b742][m742];
        end
    endgenerate
    generate 
        localparam integer b743 = 15;
        for (m743 = 0; m743 < 16; m743 = m743 + 1) 
        begin: inbit743
            assign data_11[m743 + b743*16 + a26*28*16] = data_11_array[a26][b743][m743];
        end
    endgenerate
    generate 
        localparam integer b744 = 16;
        for (m744 = 0; m744 < 16; m744 = m744 + 1) 
        begin: inbit744
            assign data_11[m744 + b744*16 + a26*28*16] = data_11_array[a26][b744][m744];
        end
    endgenerate
    generate 
        localparam integer b745 = 17;
        for (m745 = 0; m745 < 16; m745 = m745 + 1) 
        begin: inbit745
            assign data_11[m745 + b745*16 + a26*28*16] = data_11_array[a26][b745][m745];
        end
    endgenerate
    generate 
        localparam integer b746 = 18;
        for (m746 = 0; m746 < 16; m746 = m746 + 1) 
        begin: inbit746
            assign data_11[m746 + b746*16 + a26*28*16] = data_11_array[a26][b746][m746];
        end
    endgenerate
    generate 
        localparam integer b747 = 19;
        for (m747 = 0; m747 < 16; m747 = m747 + 1) 
        begin: inbit747
            assign data_11[m747 + b747*16 + a26*28*16] = data_11_array[a26][b747][m747];
        end
    endgenerate
    generate 
        localparam integer b748 = 20;
        for (m748 = 0; m748 < 16; m748 = m748 + 1) 
        begin: inbit748
            assign data_11[m748 + b748*16 + a26*28*16] = data_11_array[a26][b748][m748];
        end
    endgenerate
    generate 
        localparam integer b749 = 21;
        for (m749 = 0; m749 < 16; m749 = m749 + 1) 
        begin: inbit749
            assign data_11[m749 + b749*16 + a26*28*16] = data_11_array[a26][b749][m749];
        end
    endgenerate
    generate 
        localparam integer b750 = 22;
        for (m750 = 0; m750 < 16; m750 = m750 + 1) 
        begin: inbit750
            assign data_11[m750 + b750*16 + a26*28*16] = data_11_array[a26][b750][m750];
        end
    endgenerate
    generate 
        localparam integer b751 = 23;
        for (m751 = 0; m751 < 16; m751 = m751 + 1) 
        begin: inbit751
            assign data_11[m751 + b751*16 + a26*28*16] = data_11_array[a26][b751][m751];
        end
    endgenerate
    generate 
        localparam integer b752 = 24;
        for (m752 = 0; m752 < 16; m752 = m752 + 1) 
        begin: inbit752
            assign data_11[m752 + b752*16 + a26*28*16] = data_11_array[a26][b752][m752];
        end
    endgenerate
    generate 
        localparam integer b753 = 25;
        for (m753 = 0; m753 < 16; m753 = m753 + 1) 
        begin: inbit753
            assign data_11[m753 + b753*16 + a26*28*16] = data_11_array[a26][b753][m753];
        end
    endgenerate
    generate 
        localparam integer b754 = 26;
        for (m754 = 0; m754 < 16; m754 = m754 + 1) 
        begin: inbit754
            assign data_11[m754 + b754*16 + a26*28*16] = data_11_array[a26][b754][m754];
        end
    endgenerate
    generate 
        localparam integer b755 = 27;
        for (m755 = 0; m755 < 16; m755 = m755 + 1) 
        begin: inbit755
            assign data_11[m755 + b755*16 + a26*28*16] = data_11_array[a26][b755][m755];
        end
    endgenerate
    localparam integer a27 = 27;
    generate 
        localparam integer b756 = 0;
        for (m756 = 0; m756 < 16; m756 = m756 + 1) 
        begin: inbit756
            assign data_11[m756 + b756*16 + a27*28*16] = data_11_array[a27][b756][m756];
        end
    endgenerate
    generate 
        localparam integer b757 = 1;
        for (m757 = 0; m757 < 16; m757 = m757 + 1) 
        begin: inbit757
            assign data_11[m757 + b757*16 + a27*28*16] = data_11_array[a27][b757][m757];
        end
    endgenerate
    generate 
        localparam integer b758 = 2;
        for (m758 = 0; m758 < 16; m758 = m758 + 1) 
        begin: inbit758
            assign data_11[m758 + b758*16 + a27*28*16] = data_11_array[a27][b758][m758];
        end
    endgenerate
    generate 
        localparam integer b759 = 3;
        for (m759 = 0; m759 < 16; m759 = m759 + 1) 
        begin: inbit759
            assign data_11[m759 + b759*16 + a27*28*16] = data_11_array[a27][b759][m759];
        end
    endgenerate
    generate 
        localparam integer b760 = 4;
        for (m760 = 0; m760 < 16; m760 = m760 + 1) 
        begin: inbit760
            assign data_11[m760 + b760*16 + a27*28*16] = data_11_array[a27][b760][m760];
        end
    endgenerate
    generate 
        localparam integer b761 = 5;
        for (m761 = 0; m761 < 16; m761 = m761 + 1) 
        begin: inbit761
            assign data_11[m761 + b761*16 + a27*28*16] = data_11_array[a27][b761][m761];
        end
    endgenerate
    generate 
        localparam integer b762 = 6;
        for (m762 = 0; m762 < 16; m762 = m762 + 1) 
        begin: inbit762
            assign data_11[m762 + b762*16 + a27*28*16] = data_11_array[a27][b762][m762];
        end
    endgenerate
    generate 
        localparam integer b763 = 7;
        for (m763 = 0; m763 < 16; m763 = m763 + 1) 
        begin: inbit763
            assign data_11[m763 + b763*16 + a27*28*16] = data_11_array[a27][b763][m763];
        end
    endgenerate
    generate 
        localparam integer b764 = 8;
        for (m764 = 0; m764 < 16; m764 = m764 + 1) 
        begin: inbit764
            assign data_11[m764 + b764*16 + a27*28*16] = data_11_array[a27][b764][m764];
        end
    endgenerate
    generate 
        localparam integer b765 = 9;
        for (m765 = 0; m765 < 16; m765 = m765 + 1) 
        begin: inbit765
            assign data_11[m765 + b765*16 + a27*28*16] = data_11_array[a27][b765][m765];
        end
    endgenerate
    generate 
        localparam integer b766 = 10;
        for (m766 = 0; m766 < 16; m766 = m766 + 1) 
        begin: inbit766
            assign data_11[m766 + b766*16 + a27*28*16] = data_11_array[a27][b766][m766];
        end
    endgenerate
    generate 
        localparam integer b767 = 11;
        for (m767 = 0; m767 < 16; m767 = m767 + 1) 
        begin: inbit767
            assign data_11[m767 + b767*16 + a27*28*16] = data_11_array[a27][b767][m767];
        end
    endgenerate
    generate 
        localparam integer b768 = 12;
        for (m768 = 0; m768 < 16; m768 = m768 + 1) 
        begin: inbit768
            assign data_11[m768 + b768*16 + a27*28*16] = data_11_array[a27][b768][m768];
        end
    endgenerate
    generate 
        localparam integer b769 = 13;
        for (m769 = 0; m769 < 16; m769 = m769 + 1) 
        begin: inbit769
            assign data_11[m769 + b769*16 + a27*28*16] = data_11_array[a27][b769][m769];
        end
    endgenerate
    generate 
        localparam integer b770 = 14;
        for (m770 = 0; m770 < 16; m770 = m770 + 1) 
        begin: inbit770
            assign data_11[m770 + b770*16 + a27*28*16] = data_11_array[a27][b770][m770];
        end
    endgenerate
    generate 
        localparam integer b771 = 15;
        for (m771 = 0; m771 < 16; m771 = m771 + 1) 
        begin: inbit771
            assign data_11[m771 + b771*16 + a27*28*16] = data_11_array[a27][b771][m771];
        end
    endgenerate
    generate 
        localparam integer b772 = 16;
        for (m772 = 0; m772 < 16; m772 = m772 + 1) 
        begin: inbit772
            assign data_11[m772 + b772*16 + a27*28*16] = data_11_array[a27][b772][m772];
        end
    endgenerate
    generate 
        localparam integer b773 = 17;
        for (m773 = 0; m773 < 16; m773 = m773 + 1) 
        begin: inbit773
            assign data_11[m773 + b773*16 + a27*28*16] = data_11_array[a27][b773][m773];
        end
    endgenerate
    generate 
        localparam integer b774 = 18;
        for (m774 = 0; m774 < 16; m774 = m774 + 1) 
        begin: inbit774
            assign data_11[m774 + b774*16 + a27*28*16] = data_11_array[a27][b774][m774];
        end
    endgenerate
    generate 
        localparam integer b775 = 19;
        for (m775 = 0; m775 < 16; m775 = m775 + 1) 
        begin: inbit775
            assign data_11[m775 + b775*16 + a27*28*16] = data_11_array[a27][b775][m775];
        end
    endgenerate
    generate 
        localparam integer b776 = 20;
        for (m776 = 0; m776 < 16; m776 = m776 + 1) 
        begin: inbit776
            assign data_11[m776 + b776*16 + a27*28*16] = data_11_array[a27][b776][m776];
        end
    endgenerate
    generate 
        localparam integer b777 = 21;
        for (m777 = 0; m777 < 16; m777 = m777 + 1) 
        begin: inbit777
            assign data_11[m777 + b777*16 + a27*28*16] = data_11_array[a27][b777][m777];
        end
    endgenerate
    generate 
        localparam integer b778 = 22;
        for (m778 = 0; m778 < 16; m778 = m778 + 1) 
        begin: inbit778
            assign data_11[m778 + b778*16 + a27*28*16] = data_11_array[a27][b778][m778];
        end
    endgenerate
    generate 
        localparam integer b779 = 23;
        for (m779 = 0; m779 < 16; m779 = m779 + 1) 
        begin: inbit779
            assign data_11[m779 + b779*16 + a27*28*16] = data_11_array[a27][b779][m779];
        end
    endgenerate
    generate 
        localparam integer b780 = 24;
        for (m780 = 0; m780 < 16; m780 = m780 + 1) 
        begin: inbit780
            assign data_11[m780 + b780*16 + a27*28*16] = data_11_array[a27][b780][m780];
        end
    endgenerate
    generate 
        localparam integer b781 = 25;
        for (m781 = 0; m781 < 16; m781 = m781 + 1) 
        begin: inbit781
            assign data_11[m781 + b781*16 + a27*28*16] = data_11_array[a27][b781][m781];
        end
    endgenerate
    generate 
        localparam integer b782 = 26;
        for (m782 = 0; m782 < 16; m782 = m782 + 1) 
        begin: inbit782
            assign data_11[m782 + b782*16 + a27*28*16] = data_11_array[a27][b782][m782];
        end
    endgenerate
    generate 
        localparam integer b783 = 27;
        for (m783 = 0; m783 < 16; m783 = m783 + 1) 
        begin: inbit783
            assign data_11[m783 + b783*16 + a27*28*16] = data_11_array[a27][b783][m783];
        end
    endgenerate

  
  
  ////ROW 0
  generate
    localparam integer j0 = 0;
    for (i0 = 0; i0 < 24; i0 = i0 + 1)
    begin: addbit0
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j0+0][i0+0]), .Out(multi0[0][i0]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j0+0][i0+1]), .Out(multi0[1][i0]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j0+0][i0+2]), .Out(multi0[2][i0]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j0+0][i0+3]), .Out(multi0[3][i0]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j0+0][i0+4]), .Out(multi0[4][i0]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j0+1][i0+0]), .Out(multi0[5][i0]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j0+1][i0+1]), .Out(multi0[6][i0]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j0+1][i0+2]), .Out(multi0[7][i0]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j0+1][i0+3]), .Out(multi0[8][i0]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j0+1][i0+4]), .Out(multi0[9][i0]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j0+2][i0+0]), .Out(multi0[10][i0]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j0+2][i0+1]), .Out(multi0[11][i0]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j0+2][i0+2]), .Out(multi0[12][i0]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j0+2][i0+3]), .Out(multi0[13][i0]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j0+2][i0+4]), .Out(multi0[14][i0]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j0+3][i0+0]), .Out(multi0[15][i0]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j0+3][i0+1]), .Out(multi0[16][i0]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j0+3][i0+2]), .Out(multi0[17][i0]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j0+3][i0+3]), .Out(multi0[18][i0]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j0+3][i0+4]), .Out(multi0[19][i0]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j0+4][i0+0]), .Out(multi0[20][i0]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j0+4][i0+1]), .Out(multi0[21][i0]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j0+4][i0+2]), .Out(multi0[22][i0]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j0+4][i0+3]), .Out(multi0[23][i0]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j0+4][i0+4]), .Out(multi0[24][i0]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi0[0][i0]), .B(multi0[1][i0]), .Out(sum0[0][i0]));
      FP16_Add stage026(.A(multi0[2][i0]), .B(multi0[3][i0]), .Out(sum0[1][i0]));
      FP16_Add stage027(.A(multi0[4][i0]), .B(multi0[5][i0]), .Out(sum0[2][i0]));
      FP16_Add stage028(.A(multi0[6][i0]), .B(multi0[7][i0]), .Out(sum0[3][i0]));
      FP16_Add stage029(.A(multi0[8][i0]), .B(multi0[9][i0]), .Out(sum0[4][i0]));
      FP16_Add stage030(.A(multi0[10][i0]), .B(multi0[11][i0]), .Out(sum0[5][i0]));
      FP16_Add stage031(.A(multi0[12][i0]), .B(multi0[13][i0]), .Out(sum0[6][i0]));
      FP16_Add stage032(.A(multi0[14][i0]), .B(multi0[15][i0]), .Out(sum0[7][i0]));
      FP16_Add stage033(.A(multi0[16][i0]), .B(multi0[17][i0]), .Out(sum0[8][i0]));
      FP16_Add stage034(.A(multi0[18][i0]), .B(multi0[19][i0]), .Out(sum0[9][i0]));
      FP16_Add stage035(.A(multi0[20][i0]), .B(multi0[21][i0]), .Out(sum0[10][i0]));
      FP16_Add stage036(.A(multi0[22][i0]), .B(multi0[23][i0]), .Out(sum0[11][i0]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum0[0][i0]), .B(sum0[1][i0]), .Out(sum0[12][i0]));
      FP16_Add stage038(.A(sum0[2][i0]), .B(sum0[3][i0]), .Out(sum0[13][i0]));
      FP16_Add stage039(.A(sum0[4][i0]), .B(sum0[5][i0]), .Out(sum0[14][i0]));
      FP16_Add stage040(.A(sum0[6][i0]), .B(sum0[7][i0]), .Out(sum0[15][i0]));
      FP16_Add stage041(.A(sum0[8][i0]), .B(sum0[9][i0]), .Out(sum0[16][i0]));
      FP16_Add stage042(.A(sum0[10][i0]), .B(sum0[11][i0]), .Out(sum0[17][i0]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum0[12][i0]), .B(sum0[13][i0]), .Out(sum0[18][i0]));
      FP16_Add stage044(.A(sum0[14][i0]), .B(sum0[15][i0]), .Out(sum0[19][i0]));
      FP16_Add stage045(.A(sum0[16][i0]), .B(sum0[17][i0]), .Out(sum0[20][i0]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum0[18][i0]), .B(sum0[19][i0]), .Out(sum0[21][i0]));
      FP16_Add stage047(.A(sum0[20][i0]), .B(multi0[24][i0]), .Out(sum0[22][i0]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum0[21][i0]), .B(sum0[22][i0]), .Out(sum0[23][i0]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum0[23][i0]), .B(feature1Bias), .Out(data_11_array[j0][i0]));
    end
  endgenerate
  
  ////ROW 1
  generate
    localparam integer j1 = 1;
    for (i1 = 0; i1 < 24; i1 = i1 + 1)
    begin: addbit1
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j1+0][i1+0]), .Out(multi1[0][i1]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j1+0][i1+1]), .Out(multi1[1][i1]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j1+0][i1+2]), .Out(multi1[2][i1]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j1+0][i1+3]), .Out(multi1[3][i1]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j1+0][i1+4]), .Out(multi1[4][i1]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j1+1][i1+0]), .Out(multi1[5][i1]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j1+1][i1+1]), .Out(multi1[6][i1]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j1+1][i1+2]), .Out(multi1[7][i1]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j1+1][i1+3]), .Out(multi1[8][i1]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j1+1][i1+4]), .Out(multi1[9][i1]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j1+2][i1+0]), .Out(multi1[10][i1]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j1+2][i1+1]), .Out(multi1[11][i1]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j1+2][i1+2]), .Out(multi1[12][i1]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j1+2][i1+3]), .Out(multi1[13][i1]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j1+2][i1+4]), .Out(multi1[14][i1]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j1+3][i1+0]), .Out(multi1[15][i1]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j1+3][i1+1]), .Out(multi1[16][i1]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j1+3][i1+2]), .Out(multi1[17][i1]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j1+3][i1+3]), .Out(multi1[18][i1]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j1+3][i1+4]), .Out(multi1[19][i1]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j1+4][i1+0]), .Out(multi1[20][i1]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j1+4][i1+1]), .Out(multi1[21][i1]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j1+4][i1+2]), .Out(multi1[22][i1]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j1+4][i1+3]), .Out(multi1[23][i1]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j1+4][i1+4]), .Out(multi1[24][i1]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi1[0][i1]), .B(multi1[1][i1]), .Out(sum1[0][i1]));
      FP16_Add stage026(.A(multi1[2][i1]), .B(multi1[3][i1]), .Out(sum1[1][i1]));
      FP16_Add stage027(.A(multi1[4][i1]), .B(multi1[5][i1]), .Out(sum1[2][i1]));
      FP16_Add stage028(.A(multi1[6][i1]), .B(multi1[7][i1]), .Out(sum1[3][i1]));
      FP16_Add stage029(.A(multi1[8][i1]), .B(multi1[9][i1]), .Out(sum1[4][i1]));
      FP16_Add stage030(.A(multi1[10][i1]), .B(multi1[11][i1]), .Out(sum1[5][i1]));
      FP16_Add stage031(.A(multi1[12][i1]), .B(multi1[13][i1]), .Out(sum1[6][i1]));
      FP16_Add stage032(.A(multi1[14][i1]), .B(multi1[15][i1]), .Out(sum1[7][i1]));
      FP16_Add stage033(.A(multi1[16][i1]), .B(multi1[17][i1]), .Out(sum1[8][i1]));
      FP16_Add stage034(.A(multi1[18][i1]), .B(multi1[19][i1]), .Out(sum1[9][i1]));
      FP16_Add stage035(.A(multi1[20][i1]), .B(multi1[21][i1]), .Out(sum1[10][i1]));
      FP16_Add stage036(.A(multi1[22][i1]), .B(multi1[23][i1]), .Out(sum1[11][i1]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum1[0][i1]), .B(sum1[1][i1]), .Out(sum1[12][i1]));
      FP16_Add stage038(.A(sum1[2][i1]), .B(sum1[3][i1]), .Out(sum1[13][i1]));
      FP16_Add stage039(.A(sum1[4][i1]), .B(sum1[5][i1]), .Out(sum1[14][i1]));
      FP16_Add stage040(.A(sum1[6][i1]), .B(sum1[7][i1]), .Out(sum1[15][i1]));
      FP16_Add stage041(.A(sum1[8][i1]), .B(sum1[9][i1]), .Out(sum1[16][i1]));
      FP16_Add stage042(.A(sum1[10][i1]), .B(sum1[11][i1]), .Out(sum1[17][i1]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum1[12][i1]), .B(sum1[13][i1]), .Out(sum1[18][i1]));
      FP16_Add stage044(.A(sum1[14][i1]), .B(sum1[15][i1]), .Out(sum1[19][i1]));
      FP16_Add stage045(.A(sum1[16][i1]), .B(sum1[17][i1]), .Out(sum1[20][i1]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum1[18][i1]), .B(sum1[19][i1]), .Out(sum1[21][i1]));
      FP16_Add stage047(.A(sum1[20][i1]), .B(multi1[24][i1]), .Out(sum1[22][i1]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum1[21][i1]), .B(sum1[22][i1]), .Out(sum1[23][i1]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum1[23][i1]), .B(feature1Bias), .Out(data_11_array[j1][i1]));
    end
  endgenerate
  
  ////ROW 2
  generate
    localparam integer j2 = 2;
    for (i2 = 0; i2 < 24; i2 = i2 + 1)
    begin: addbit2
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j2+0][i2+0]), .Out(multi2[0][i2]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j2+0][i2+1]), .Out(multi2[1][i2]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j2+0][i2+2]), .Out(multi2[2][i2]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j2+0][i2+3]), .Out(multi2[3][i2]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j2+0][i2+4]), .Out(multi2[4][i2]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j2+1][i2+0]), .Out(multi2[5][i2]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j2+1][i2+1]), .Out(multi2[6][i2]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j2+1][i2+2]), .Out(multi2[7][i2]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j2+1][i2+3]), .Out(multi2[8][i2]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j2+1][i2+4]), .Out(multi2[9][i2]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j2+2][i2+0]), .Out(multi2[10][i2]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j2+2][i2+1]), .Out(multi2[11][i2]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j2+2][i2+2]), .Out(multi2[12][i2]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j2+2][i2+3]), .Out(multi2[13][i2]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j2+2][i2+4]), .Out(multi2[14][i2]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j2+3][i2+0]), .Out(multi2[15][i2]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j2+3][i2+1]), .Out(multi2[16][i2]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j2+3][i2+2]), .Out(multi2[17][i2]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j2+3][i2+3]), .Out(multi2[18][i2]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j2+3][i2+4]), .Out(multi2[19][i2]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j2+4][i2+0]), .Out(multi2[20][i2]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j2+4][i2+1]), .Out(multi2[21][i2]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j2+4][i2+2]), .Out(multi2[22][i2]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j2+4][i2+3]), .Out(multi2[23][i2]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j2+4][i2+4]), .Out(multi2[24][i2]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi2[0][i2]), .B(multi2[1][i2]), .Out(sum2[0][i2]));
      FP16_Add stage026(.A(multi2[2][i2]), .B(multi2[3][i2]), .Out(sum2[1][i2]));
      FP16_Add stage027(.A(multi2[4][i2]), .B(multi2[5][i2]), .Out(sum2[2][i2]));
      FP16_Add stage028(.A(multi2[6][i2]), .B(multi2[7][i2]), .Out(sum2[3][i2]));
      FP16_Add stage029(.A(multi2[8][i2]), .B(multi2[9][i2]), .Out(sum2[4][i2]));
      FP16_Add stage030(.A(multi2[10][i2]), .B(multi2[11][i2]), .Out(sum2[5][i2]));
      FP16_Add stage031(.A(multi2[12][i2]), .B(multi2[13][i2]), .Out(sum2[6][i2]));
      FP16_Add stage032(.A(multi2[14][i2]), .B(multi2[15][i2]), .Out(sum2[7][i2]));
      FP16_Add stage033(.A(multi2[16][i2]), .B(multi2[17][i2]), .Out(sum2[8][i2]));
      FP16_Add stage034(.A(multi2[18][i2]), .B(multi2[19][i2]), .Out(sum2[9][i2]));
      FP16_Add stage035(.A(multi2[20][i2]), .B(multi2[21][i2]), .Out(sum2[10][i2]));
      FP16_Add stage036(.A(multi2[22][i2]), .B(multi2[23][i2]), .Out(sum2[11][i2]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum2[0][i2]), .B(sum2[1][i2]), .Out(sum2[12][i2]));
      FP16_Add stage038(.A(sum2[2][i2]), .B(sum2[3][i2]), .Out(sum2[13][i2]));
      FP16_Add stage039(.A(sum2[4][i2]), .B(sum2[5][i2]), .Out(sum2[14][i2]));
      FP16_Add stage040(.A(sum2[6][i2]), .B(sum2[7][i2]), .Out(sum2[15][i2]));
      FP16_Add stage041(.A(sum2[8][i2]), .B(sum2[9][i2]), .Out(sum2[16][i2]));
      FP16_Add stage042(.A(sum2[10][i2]), .B(sum2[11][i2]), .Out(sum2[17][i2]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum2[12][i2]), .B(sum2[13][i2]), .Out(sum2[18][i2]));
      FP16_Add stage044(.A(sum2[14][i2]), .B(sum2[15][i2]), .Out(sum2[19][i2]));
      FP16_Add stage045(.A(sum2[16][i2]), .B(sum2[17][i2]), .Out(sum2[20][i2]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum2[18][i2]), .B(sum2[19][i2]), .Out(sum2[21][i2]));
      FP16_Add stage047(.A(sum2[20][i2]), .B(multi2[24][i2]), .Out(sum2[22][i2]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum2[21][i2]), .B(sum2[22][i2]), .Out(sum2[23][i2]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum2[23][i2]), .B(feature1Bias), .Out(data_11_array[j2][i2]));
    end
  endgenerate
  
  ////ROW 3
  generate
    localparam integer j3 = 3;
    for (i3 = 0; i3 < 24; i3 = i3 + 1)
    begin: addbit3
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j3+0][i3+0]), .Out(multi3[0][i3]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j3+0][i3+1]), .Out(multi3[1][i3]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j3+0][i3+2]), .Out(multi3[2][i3]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j3+0][i3+3]), .Out(multi3[3][i3]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j3+0][i3+4]), .Out(multi3[4][i3]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j3+1][i3+0]), .Out(multi3[5][i3]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j3+1][i3+1]), .Out(multi3[6][i3]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j3+1][i3+2]), .Out(multi3[7][i3]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j3+1][i3+3]), .Out(multi3[8][i3]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j3+1][i3+4]), .Out(multi3[9][i3]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j3+2][i3+0]), .Out(multi3[10][i3]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j3+2][i3+1]), .Out(multi3[11][i3]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j3+2][i3+2]), .Out(multi3[12][i3]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j3+2][i3+3]), .Out(multi3[13][i3]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j3+2][i3+4]), .Out(multi3[14][i3]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j3+3][i3+0]), .Out(multi3[15][i3]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j3+3][i3+1]), .Out(multi3[16][i3]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j3+3][i3+2]), .Out(multi3[17][i3]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j3+3][i3+3]), .Out(multi3[18][i3]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j3+3][i3+4]), .Out(multi3[19][i3]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j3+4][i3+0]), .Out(multi3[20][i3]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j3+4][i3+1]), .Out(multi3[21][i3]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j3+4][i3+2]), .Out(multi3[22][i3]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j3+4][i3+3]), .Out(multi3[23][i3]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j3+4][i3+4]), .Out(multi3[24][i3]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi3[0][i3]), .B(multi3[1][i3]), .Out(sum3[0][i3]));
      FP16_Add stage026(.A(multi3[2][i3]), .B(multi3[3][i3]), .Out(sum3[1][i3]));
      FP16_Add stage027(.A(multi3[4][i3]), .B(multi3[5][i3]), .Out(sum3[2][i3]));
      FP16_Add stage028(.A(multi3[6][i3]), .B(multi3[7][i3]), .Out(sum3[3][i3]));
      FP16_Add stage029(.A(multi3[8][i3]), .B(multi3[9][i3]), .Out(sum3[4][i3]));
      FP16_Add stage030(.A(multi3[10][i3]), .B(multi3[11][i3]), .Out(sum3[5][i3]));
      FP16_Add stage031(.A(multi3[12][i3]), .B(multi3[13][i3]), .Out(sum3[6][i3]));
      FP16_Add stage032(.A(multi3[14][i3]), .B(multi3[15][i3]), .Out(sum3[7][i3]));
      FP16_Add stage033(.A(multi3[16][i3]), .B(multi3[17][i3]), .Out(sum3[8][i3]));
      FP16_Add stage034(.A(multi3[18][i3]), .B(multi3[19][i3]), .Out(sum3[9][i3]));
      FP16_Add stage035(.A(multi3[20][i3]), .B(multi3[21][i3]), .Out(sum3[10][i3]));
      FP16_Add stage036(.A(multi3[22][i3]), .B(multi3[23][i3]), .Out(sum3[11][i3]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum3[0][i3]), .B(sum3[1][i3]), .Out(sum3[12][i3]));
      FP16_Add stage038(.A(sum3[2][i3]), .B(sum3[3][i3]), .Out(sum3[13][i3]));
      FP16_Add stage039(.A(sum3[4][i3]), .B(sum3[5][i3]), .Out(sum3[14][i3]));
      FP16_Add stage040(.A(sum3[6][i3]), .B(sum3[7][i3]), .Out(sum3[15][i3]));
      FP16_Add stage041(.A(sum3[8][i3]), .B(sum3[9][i3]), .Out(sum3[16][i3]));
      FP16_Add stage042(.A(sum3[10][i3]), .B(sum3[11][i3]), .Out(sum3[17][i3]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum3[12][i3]), .B(sum3[13][i3]), .Out(sum3[18][i3]));
      FP16_Add stage044(.A(sum3[14][i3]), .B(sum3[15][i3]), .Out(sum3[19][i3]));
      FP16_Add stage045(.A(sum3[16][i3]), .B(sum3[17][i3]), .Out(sum3[20][i3]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum3[18][i3]), .B(sum3[19][i3]), .Out(sum3[21][i3]));
      FP16_Add stage047(.A(sum3[20][i3]), .B(multi3[24][i3]), .Out(sum3[22][i3]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum3[21][i3]), .B(sum3[22][i3]), .Out(sum3[23][i3]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum3[23][i3]), .B(feature1Bias), .Out(data_11_array[j3][i3]));
    end
  endgenerate
  
  ////ROW 4
  generate
    localparam integer j4 = 4;
    for (i4 = 0; i4 < 24; i4 = i4 + 1)
    begin: addbit4
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j4+0][i4+0]), .Out(multi4[0][i4]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j4+0][i4+1]), .Out(multi4[1][i4]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j4+0][i4+2]), .Out(multi4[2][i4]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j4+0][i4+3]), .Out(multi4[3][i4]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j4+0][i4+4]), .Out(multi4[4][i4]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j4+1][i4+0]), .Out(multi4[5][i4]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j4+1][i4+1]), .Out(multi4[6][i4]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j4+1][i4+2]), .Out(multi4[7][i4]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j4+1][i4+3]), .Out(multi4[8][i4]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j4+1][i4+4]), .Out(multi4[9][i4]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j4+2][i4+0]), .Out(multi4[10][i4]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j4+2][i4+1]), .Out(multi4[11][i4]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j4+2][i4+2]), .Out(multi4[12][i4]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j4+2][i4+3]), .Out(multi4[13][i4]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j4+2][i4+4]), .Out(multi4[14][i4]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j4+3][i4+0]), .Out(multi4[15][i4]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j4+3][i4+1]), .Out(multi4[16][i4]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j4+3][i4+2]), .Out(multi4[17][i4]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j4+3][i4+3]), .Out(multi4[18][i4]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j4+3][i4+4]), .Out(multi4[19][i4]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j4+4][i4+0]), .Out(multi4[20][i4]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j4+4][i4+1]), .Out(multi4[21][i4]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j4+4][i4+2]), .Out(multi4[22][i4]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j4+4][i4+3]), .Out(multi4[23][i4]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j4+4][i4+4]), .Out(multi4[24][i4]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi4[0][i4]), .B(multi4[1][i4]), .Out(sum4[0][i4]));
      FP16_Add stage026(.A(multi4[2][i4]), .B(multi4[3][i4]), .Out(sum4[1][i4]));
      FP16_Add stage027(.A(multi4[4][i4]), .B(multi4[5][i4]), .Out(sum4[2][i4]));
      FP16_Add stage028(.A(multi4[6][i4]), .B(multi4[7][i4]), .Out(sum4[3][i4]));
      FP16_Add stage029(.A(multi4[8][i4]), .B(multi4[9][i4]), .Out(sum4[4][i4]));
      FP16_Add stage030(.A(multi4[10][i4]), .B(multi4[11][i4]), .Out(sum4[5][i4]));
      FP16_Add stage031(.A(multi4[12][i4]), .B(multi4[13][i4]), .Out(sum4[6][i4]));
      FP16_Add stage032(.A(multi4[14][i4]), .B(multi4[15][i4]), .Out(sum4[7][i4]));
      FP16_Add stage033(.A(multi4[16][i4]), .B(multi4[17][i4]), .Out(sum4[8][i4]));
      FP16_Add stage034(.A(multi4[18][i4]), .B(multi4[19][i4]), .Out(sum4[9][i4]));
      FP16_Add stage035(.A(multi4[20][i4]), .B(multi4[21][i4]), .Out(sum4[10][i4]));
      FP16_Add stage036(.A(multi4[22][i4]), .B(multi4[23][i4]), .Out(sum4[11][i4]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum4[0][i4]), .B(sum4[1][i4]), .Out(sum4[12][i4]));
      FP16_Add stage038(.A(sum4[2][i4]), .B(sum4[3][i4]), .Out(sum4[13][i4]));
      FP16_Add stage039(.A(sum4[4][i4]), .B(sum4[5][i4]), .Out(sum4[14][i4]));
      FP16_Add stage040(.A(sum4[6][i4]), .B(sum4[7][i4]), .Out(sum4[15][i4]));
      FP16_Add stage041(.A(sum4[8][i4]), .B(sum4[9][i4]), .Out(sum4[16][i4]));
      FP16_Add stage042(.A(sum4[10][i4]), .B(sum4[11][i4]), .Out(sum4[17][i4]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum4[12][i4]), .B(sum4[13][i4]), .Out(sum4[18][i4]));
      FP16_Add stage044(.A(sum4[14][i4]), .B(sum4[15][i4]), .Out(sum4[19][i4]));
      FP16_Add stage045(.A(sum4[16][i4]), .B(sum4[17][i4]), .Out(sum4[20][i4]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum4[18][i4]), .B(sum4[19][i4]), .Out(sum4[21][i4]));
      FP16_Add stage047(.A(sum4[20][i4]), .B(multi4[24][i4]), .Out(sum4[22][i4]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum4[21][i4]), .B(sum4[22][i4]), .Out(sum4[23][i4]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum4[23][i4]), .B(feature1Bias), .Out(data_11_array[j4][i4]));
    end
  endgenerate
  
  ////ROW 5
  generate
    localparam integer j5 = 5;
    for (i5 = 0; i5 < 24; i5 = i5 + 1)
    begin: addbit5
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j5+0][i5+0]), .Out(multi5[0][i5]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j5+0][i5+1]), .Out(multi5[1][i5]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j5+0][i5+2]), .Out(multi5[2][i5]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j5+0][i5+3]), .Out(multi5[3][i5]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j5+0][i5+4]), .Out(multi5[4][i5]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j5+1][i5+0]), .Out(multi5[5][i5]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j5+1][i5+1]), .Out(multi5[6][i5]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j5+1][i5+2]), .Out(multi5[7][i5]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j5+1][i5+3]), .Out(multi5[8][i5]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j5+1][i5+4]), .Out(multi5[9][i5]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j5+2][i5+0]), .Out(multi5[10][i5]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j5+2][i5+1]), .Out(multi5[11][i5]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j5+2][i5+2]), .Out(multi5[12][i5]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j5+2][i5+3]), .Out(multi5[13][i5]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j5+2][i5+4]), .Out(multi5[14][i5]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j5+3][i5+0]), .Out(multi5[15][i5]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j5+3][i5+1]), .Out(multi5[16][i5]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j5+3][i5+2]), .Out(multi5[17][i5]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j5+3][i5+3]), .Out(multi5[18][i5]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j5+3][i5+4]), .Out(multi5[19][i5]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j5+4][i5+0]), .Out(multi5[20][i5]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j5+4][i5+1]), .Out(multi5[21][i5]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j5+4][i5+2]), .Out(multi5[22][i5]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j5+4][i5+3]), .Out(multi5[23][i5]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j5+4][i5+4]), .Out(multi5[24][i5]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi5[0][i5]), .B(multi5[1][i5]), .Out(sum5[0][i5]));
      FP16_Add stage026(.A(multi5[2][i5]), .B(multi5[3][i5]), .Out(sum5[1][i5]));
      FP16_Add stage027(.A(multi5[4][i5]), .B(multi5[5][i5]), .Out(sum5[2][i5]));
      FP16_Add stage028(.A(multi5[6][i5]), .B(multi5[7][i5]), .Out(sum5[3][i5]));
      FP16_Add stage029(.A(multi5[8][i5]), .B(multi5[9][i5]), .Out(sum5[4][i5]));
      FP16_Add stage030(.A(multi5[10][i5]), .B(multi5[11][i5]), .Out(sum5[5][i5]));
      FP16_Add stage031(.A(multi5[12][i5]), .B(multi5[13][i5]), .Out(sum5[6][i5]));
      FP16_Add stage032(.A(multi5[14][i5]), .B(multi5[15][i5]), .Out(sum5[7][i5]));
      FP16_Add stage033(.A(multi5[16][i5]), .B(multi5[17][i5]), .Out(sum5[8][i5]));
      FP16_Add stage034(.A(multi5[18][i5]), .B(multi5[19][i5]), .Out(sum5[9][i5]));
      FP16_Add stage035(.A(multi5[20][i5]), .B(multi5[21][i5]), .Out(sum5[10][i5]));
      FP16_Add stage036(.A(multi5[22][i5]), .B(multi5[23][i5]), .Out(sum5[11][i5]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum5[0][i5]), .B(sum5[1][i5]), .Out(sum5[12][i5]));
      FP16_Add stage038(.A(sum5[2][i5]), .B(sum5[3][i5]), .Out(sum5[13][i5]));
      FP16_Add stage039(.A(sum5[4][i5]), .B(sum5[5][i5]), .Out(sum5[14][i5]));
      FP16_Add stage040(.A(sum5[6][i5]), .B(sum5[7][i5]), .Out(sum5[15][i5]));
      FP16_Add stage041(.A(sum5[8][i5]), .B(sum5[9][i5]), .Out(sum5[16][i5]));
      FP16_Add stage042(.A(sum5[10][i5]), .B(sum5[11][i5]), .Out(sum5[17][i5]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum5[12][i5]), .B(sum5[13][i5]), .Out(sum5[18][i5]));
      FP16_Add stage044(.A(sum5[14][i5]), .B(sum5[15][i5]), .Out(sum5[19][i5]));
      FP16_Add stage045(.A(sum5[16][i5]), .B(sum5[17][i5]), .Out(sum5[20][i5]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum5[18][i5]), .B(sum5[19][i5]), .Out(sum5[21][i5]));
      FP16_Add stage047(.A(sum5[20][i5]), .B(multi5[24][i5]), .Out(sum5[22][i5]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum5[21][i5]), .B(sum5[22][i5]), .Out(sum5[23][i5]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum5[23][i5]), .B(feature1Bias), .Out(data_11_array[j5][i5]));
    end
  endgenerate
  
  ////ROW 6
  generate
    localparam integer j6 = 6;
    for (i6 = 0; i6 < 24; i6 = i6 + 1)
    begin: addbit6
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j6+0][i6+0]), .Out(multi6[0][i6]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j6+0][i6+1]), .Out(multi6[1][i6]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j6+0][i6+2]), .Out(multi6[2][i6]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j6+0][i6+3]), .Out(multi6[3][i6]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j6+0][i6+4]), .Out(multi6[4][i6]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j6+1][i6+0]), .Out(multi6[5][i6]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j6+1][i6+1]), .Out(multi6[6][i6]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j6+1][i6+2]), .Out(multi6[7][i6]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j6+1][i6+3]), .Out(multi6[8][i6]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j6+1][i6+4]), .Out(multi6[9][i6]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j6+2][i6+0]), .Out(multi6[10][i6]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j6+2][i6+1]), .Out(multi6[11][i6]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j6+2][i6+2]), .Out(multi6[12][i6]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j6+2][i6+3]), .Out(multi6[13][i6]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j6+2][i6+4]), .Out(multi6[14][i6]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j6+3][i6+0]), .Out(multi6[15][i6]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j6+3][i6+1]), .Out(multi6[16][i6]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j6+3][i6+2]), .Out(multi6[17][i6]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j6+3][i6+3]), .Out(multi6[18][i6]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j6+3][i6+4]), .Out(multi6[19][i6]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j6+4][i6+0]), .Out(multi6[20][i6]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j6+4][i6+1]), .Out(multi6[21][i6]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j6+4][i6+2]), .Out(multi6[22][i6]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j6+4][i6+3]), .Out(multi6[23][i6]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j6+4][i6+4]), .Out(multi6[24][i6]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi6[0][i6]), .B(multi6[1][i6]), .Out(sum6[0][i6]));
      FP16_Add stage026(.A(multi6[2][i6]), .B(multi6[3][i6]), .Out(sum6[1][i6]));
      FP16_Add stage027(.A(multi6[4][i6]), .B(multi6[5][i6]), .Out(sum6[2][i6]));
      FP16_Add stage028(.A(multi6[6][i6]), .B(multi6[7][i6]), .Out(sum6[3][i6]));
      FP16_Add stage029(.A(multi6[8][i6]), .B(multi6[9][i6]), .Out(sum6[4][i6]));
      FP16_Add stage030(.A(multi6[10][i6]), .B(multi6[11][i6]), .Out(sum6[5][i6]));
      FP16_Add stage031(.A(multi6[12][i6]), .B(multi6[13][i6]), .Out(sum6[6][i6]));
      FP16_Add stage032(.A(multi6[14][i6]), .B(multi6[15][i6]), .Out(sum6[7][i6]));
      FP16_Add stage033(.A(multi6[16][i6]), .B(multi6[17][i6]), .Out(sum6[8][i6]));
      FP16_Add stage034(.A(multi6[18][i6]), .B(multi6[19][i6]), .Out(sum6[9][i6]));
      FP16_Add stage035(.A(multi6[20][i6]), .B(multi6[21][i6]), .Out(sum6[10][i6]));
      FP16_Add stage036(.A(multi6[22][i6]), .B(multi6[23][i6]), .Out(sum6[11][i6]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum6[0][i6]), .B(sum6[1][i6]), .Out(sum6[12][i6]));
      FP16_Add stage038(.A(sum6[2][i6]), .B(sum6[3][i6]), .Out(sum6[13][i6]));
      FP16_Add stage039(.A(sum6[4][i6]), .B(sum6[5][i6]), .Out(sum6[14][i6]));
      FP16_Add stage040(.A(sum6[6][i6]), .B(sum6[7][i6]), .Out(sum6[15][i6]));
      FP16_Add stage041(.A(sum6[8][i6]), .B(sum6[9][i6]), .Out(sum6[16][i6]));
      FP16_Add stage042(.A(sum6[10][i6]), .B(sum6[11][i6]), .Out(sum6[17][i6]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum6[12][i6]), .B(sum6[13][i6]), .Out(sum6[18][i6]));
      FP16_Add stage044(.A(sum6[14][i6]), .B(sum6[15][i6]), .Out(sum6[19][i6]));
      FP16_Add stage045(.A(sum6[16][i6]), .B(sum6[17][i6]), .Out(sum6[20][i6]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum6[18][i6]), .B(sum6[19][i6]), .Out(sum6[21][i6]));
      FP16_Add stage047(.A(sum6[20][i6]), .B(multi6[24][i6]), .Out(sum6[22][i6]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum6[21][i6]), .B(sum6[22][i6]), .Out(sum6[23][i6]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum6[23][i6]), .B(feature1Bias), .Out(data_11_array[j6][i6]));
    end
  endgenerate
  
  ////ROW 7
  generate
    localparam integer j7 = 7;
    for (i7 = 0; i7 < 24; i7 = i7 + 1)
    begin: addbit7
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j7+0][i7+0]), .Out(multi7[0][i7]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j7+0][i7+1]), .Out(multi7[1][i7]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j7+0][i7+2]), .Out(multi7[2][i7]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j7+0][i7+3]), .Out(multi7[3][i7]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j7+0][i7+4]), .Out(multi7[4][i7]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j7+1][i7+0]), .Out(multi7[5][i7]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j7+1][i7+1]), .Out(multi7[6][i7]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j7+1][i7+2]), .Out(multi7[7][i7]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j7+1][i7+3]), .Out(multi7[8][i7]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j7+1][i7+4]), .Out(multi7[9][i7]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j7+2][i7+0]), .Out(multi7[10][i7]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j7+2][i7+1]), .Out(multi7[11][i7]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j7+2][i7+2]), .Out(multi7[12][i7]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j7+2][i7+3]), .Out(multi7[13][i7]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j7+2][i7+4]), .Out(multi7[14][i7]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j7+3][i7+0]), .Out(multi7[15][i7]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j7+3][i7+1]), .Out(multi7[16][i7]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j7+3][i7+2]), .Out(multi7[17][i7]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j7+3][i7+3]), .Out(multi7[18][i7]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j7+3][i7+4]), .Out(multi7[19][i7]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j7+4][i7+0]), .Out(multi7[20][i7]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j7+4][i7+1]), .Out(multi7[21][i7]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j7+4][i7+2]), .Out(multi7[22][i7]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j7+4][i7+3]), .Out(multi7[23][i7]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j7+4][i7+4]), .Out(multi7[24][i7]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi7[0][i7]), .B(multi7[1][i7]), .Out(sum7[0][i7]));
      FP16_Add stage026(.A(multi7[2][i7]), .B(multi7[3][i7]), .Out(sum7[1][i7]));
      FP16_Add stage027(.A(multi7[4][i7]), .B(multi7[5][i7]), .Out(sum7[2][i7]));
      FP16_Add stage028(.A(multi7[6][i7]), .B(multi7[7][i7]), .Out(sum7[3][i7]));
      FP16_Add stage029(.A(multi7[8][i7]), .B(multi7[9][i7]), .Out(sum7[4][i7]));
      FP16_Add stage030(.A(multi7[10][i7]), .B(multi7[11][i7]), .Out(sum7[5][i7]));
      FP16_Add stage031(.A(multi7[12][i7]), .B(multi7[13][i7]), .Out(sum7[6][i7]));
      FP16_Add stage032(.A(multi7[14][i7]), .B(multi7[15][i7]), .Out(sum7[7][i7]));
      FP16_Add stage033(.A(multi7[16][i7]), .B(multi7[17][i7]), .Out(sum7[8][i7]));
      FP16_Add stage034(.A(multi7[18][i7]), .B(multi7[19][i7]), .Out(sum7[9][i7]));
      FP16_Add stage035(.A(multi7[20][i7]), .B(multi7[21][i7]), .Out(sum7[10][i7]));
      FP16_Add stage036(.A(multi7[22][i7]), .B(multi7[23][i7]), .Out(sum7[11][i7]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum7[0][i7]), .B(sum7[1][i7]), .Out(sum7[12][i7]));
      FP16_Add stage038(.A(sum7[2][i7]), .B(sum7[3][i7]), .Out(sum7[13][i7]));
      FP16_Add stage039(.A(sum7[4][i7]), .B(sum7[5][i7]), .Out(sum7[14][i7]));
      FP16_Add stage040(.A(sum7[6][i7]), .B(sum7[7][i7]), .Out(sum7[15][i7]));
      FP16_Add stage041(.A(sum7[8][i7]), .B(sum7[9][i7]), .Out(sum7[16][i7]));
      FP16_Add stage042(.A(sum7[10][i7]), .B(sum7[11][i7]), .Out(sum7[17][i7]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum7[12][i7]), .B(sum7[13][i7]), .Out(sum7[18][i7]));
      FP16_Add stage044(.A(sum7[14][i7]), .B(sum7[15][i7]), .Out(sum7[19][i7]));
      FP16_Add stage045(.A(sum7[16][i7]), .B(sum7[17][i7]), .Out(sum7[20][i7]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum7[18][i7]), .B(sum7[19][i7]), .Out(sum7[21][i7]));
      FP16_Add stage047(.A(sum7[20][i7]), .B(multi7[24][i7]), .Out(sum7[22][i7]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum7[21][i7]), .B(sum7[22][i7]), .Out(sum7[23][i7]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum7[23][i7]), .B(feature1Bias), .Out(data_11_array[j7][i7]));
    end
  endgenerate
  
  ////ROW 8
  generate
    localparam integer j8 = 8;
    for (i8 = 0; i8 < 24; i8 = i8 + 1)
    begin: addbit8
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j8+0][i8+0]), .Out(multi8[0][i8]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j8+0][i8+1]), .Out(multi8[1][i8]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j8+0][i8+2]), .Out(multi8[2][i8]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j8+0][i8+3]), .Out(multi8[3][i8]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j8+0][i8+4]), .Out(multi8[4][i8]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j8+1][i8+0]), .Out(multi8[5][i8]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j8+1][i8+1]), .Out(multi8[6][i8]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j8+1][i8+2]), .Out(multi8[7][i8]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j8+1][i8+3]), .Out(multi8[8][i8]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j8+1][i8+4]), .Out(multi8[9][i8]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j8+2][i8+0]), .Out(multi8[10][i8]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j8+2][i8+1]), .Out(multi8[11][i8]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j8+2][i8+2]), .Out(multi8[12][i8]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j8+2][i8+3]), .Out(multi8[13][i8]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j8+2][i8+4]), .Out(multi8[14][i8]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j8+3][i8+0]), .Out(multi8[15][i8]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j8+3][i8+1]), .Out(multi8[16][i8]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j8+3][i8+2]), .Out(multi8[17][i8]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j8+3][i8+3]), .Out(multi8[18][i8]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j8+3][i8+4]), .Out(multi8[19][i8]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j8+4][i8+0]), .Out(multi8[20][i8]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j8+4][i8+1]), .Out(multi8[21][i8]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j8+4][i8+2]), .Out(multi8[22][i8]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j8+4][i8+3]), .Out(multi8[23][i8]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j8+4][i8+4]), .Out(multi8[24][i8]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi8[0][i8]), .B(multi8[1][i8]), .Out(sum8[0][i8]));
      FP16_Add stage026(.A(multi8[2][i8]), .B(multi8[3][i8]), .Out(sum8[1][i8]));
      FP16_Add stage027(.A(multi8[4][i8]), .B(multi8[5][i8]), .Out(sum8[2][i8]));
      FP16_Add stage028(.A(multi8[6][i8]), .B(multi8[7][i8]), .Out(sum8[3][i8]));
      FP16_Add stage029(.A(multi8[8][i8]), .B(multi8[9][i8]), .Out(sum8[4][i8]));
      FP16_Add stage030(.A(multi8[10][i8]), .B(multi8[11][i8]), .Out(sum8[5][i8]));
      FP16_Add stage031(.A(multi8[12][i8]), .B(multi8[13][i8]), .Out(sum8[6][i8]));
      FP16_Add stage032(.A(multi8[14][i8]), .B(multi8[15][i8]), .Out(sum8[7][i8]));
      FP16_Add stage033(.A(multi8[16][i8]), .B(multi8[17][i8]), .Out(sum8[8][i8]));
      FP16_Add stage034(.A(multi8[18][i8]), .B(multi8[19][i8]), .Out(sum8[9][i8]));
      FP16_Add stage035(.A(multi8[20][i8]), .B(multi8[21][i8]), .Out(sum8[10][i8]));
      FP16_Add stage036(.A(multi8[22][i8]), .B(multi8[23][i8]), .Out(sum8[11][i8]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum8[0][i8]), .B(sum8[1][i8]), .Out(sum8[12][i8]));
      FP16_Add stage038(.A(sum8[2][i8]), .B(sum8[3][i8]), .Out(sum8[13][i8]));
      FP16_Add stage039(.A(sum8[4][i8]), .B(sum8[5][i8]), .Out(sum8[14][i8]));
      FP16_Add stage040(.A(sum8[6][i8]), .B(sum8[7][i8]), .Out(sum8[15][i8]));
      FP16_Add stage041(.A(sum8[8][i8]), .B(sum8[9][i8]), .Out(sum8[16][i8]));
      FP16_Add stage042(.A(sum8[10][i8]), .B(sum8[11][i8]), .Out(sum8[17][i8]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum8[12][i8]), .B(sum8[13][i8]), .Out(sum8[18][i8]));
      FP16_Add stage044(.A(sum8[14][i8]), .B(sum8[15][i8]), .Out(sum8[19][i8]));
      FP16_Add stage045(.A(sum8[16][i8]), .B(sum8[17][i8]), .Out(sum8[20][i8]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum8[18][i8]), .B(sum8[19][i8]), .Out(sum8[21][i8]));
      FP16_Add stage047(.A(sum8[20][i8]), .B(multi8[24][i8]), .Out(sum8[22][i8]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum8[21][i8]), .B(sum8[22][i8]), .Out(sum8[23][i8]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum8[23][i8]), .B(feature1Bias), .Out(data_11_array[j8][i8]));
    end
  endgenerate
  
  ////ROW 9
  generate
    localparam integer j9 = 9;
    for (i9 = 0; i9 < 24; i9 = i9 + 1)
    begin: addbit9
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j9+0][i9+0]), .Out(multi9[0][i9]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j9+0][i9+1]), .Out(multi9[1][i9]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j9+0][i9+2]), .Out(multi9[2][i9]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j9+0][i9+3]), .Out(multi9[3][i9]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j9+0][i9+4]), .Out(multi9[4][i9]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j9+1][i9+0]), .Out(multi9[5][i9]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j9+1][i9+1]), .Out(multi9[6][i9]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j9+1][i9+2]), .Out(multi9[7][i9]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j9+1][i9+3]), .Out(multi9[8][i9]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j9+1][i9+4]), .Out(multi9[9][i9]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j9+2][i9+0]), .Out(multi9[10][i9]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j9+2][i9+1]), .Out(multi9[11][i9]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j9+2][i9+2]), .Out(multi9[12][i9]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j9+2][i9+3]), .Out(multi9[13][i9]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j9+2][i9+4]), .Out(multi9[14][i9]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j9+3][i9+0]), .Out(multi9[15][i9]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j9+3][i9+1]), .Out(multi9[16][i9]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j9+3][i9+2]), .Out(multi9[17][i9]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j9+3][i9+3]), .Out(multi9[18][i9]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j9+3][i9+4]), .Out(multi9[19][i9]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j9+4][i9+0]), .Out(multi9[20][i9]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j9+4][i9+1]), .Out(multi9[21][i9]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j9+4][i9+2]), .Out(multi9[22][i9]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j9+4][i9+3]), .Out(multi9[23][i9]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j9+4][i9+4]), .Out(multi9[24][i9]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi9[0][i9]), .B(multi9[1][i9]), .Out(sum9[0][i9]));
      FP16_Add stage026(.A(multi9[2][i9]), .B(multi9[3][i9]), .Out(sum9[1][i9]));
      FP16_Add stage027(.A(multi9[4][i9]), .B(multi9[5][i9]), .Out(sum9[2][i9]));
      FP16_Add stage028(.A(multi9[6][i9]), .B(multi9[7][i9]), .Out(sum9[3][i9]));
      FP16_Add stage029(.A(multi9[8][i9]), .B(multi9[9][i9]), .Out(sum9[4][i9]));
      FP16_Add stage030(.A(multi9[10][i9]), .B(multi9[11][i9]), .Out(sum9[5][i9]));
      FP16_Add stage031(.A(multi9[12][i9]), .B(multi9[13][i9]), .Out(sum9[6][i9]));
      FP16_Add stage032(.A(multi9[14][i9]), .B(multi9[15][i9]), .Out(sum9[7][i9]));
      FP16_Add stage033(.A(multi9[16][i9]), .B(multi9[17][i9]), .Out(sum9[8][i9]));
      FP16_Add stage034(.A(multi9[18][i9]), .B(multi9[19][i9]), .Out(sum9[9][i9]));
      FP16_Add stage035(.A(multi9[20][i9]), .B(multi9[21][i9]), .Out(sum9[10][i9]));
      FP16_Add stage036(.A(multi9[22][i9]), .B(multi9[23][i9]), .Out(sum9[11][i9]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum9[0][i9]), .B(sum9[1][i9]), .Out(sum9[12][i9]));
      FP16_Add stage038(.A(sum9[2][i9]), .B(sum9[3][i9]), .Out(sum9[13][i9]));
      FP16_Add stage039(.A(sum9[4][i9]), .B(sum9[5][i9]), .Out(sum9[14][i9]));
      FP16_Add stage040(.A(sum9[6][i9]), .B(sum9[7][i9]), .Out(sum9[15][i9]));
      FP16_Add stage041(.A(sum9[8][i9]), .B(sum9[9][i9]), .Out(sum9[16][i9]));
      FP16_Add stage042(.A(sum9[10][i9]), .B(sum9[11][i9]), .Out(sum9[17][i9]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum9[12][i9]), .B(sum9[13][i9]), .Out(sum9[18][i9]));
      FP16_Add stage044(.A(sum9[14][i9]), .B(sum9[15][i9]), .Out(sum9[19][i9]));
      FP16_Add stage045(.A(sum9[16][i9]), .B(sum9[17][i9]), .Out(sum9[20][i9]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum9[18][i9]), .B(sum9[19][i9]), .Out(sum9[21][i9]));
      FP16_Add stage047(.A(sum9[20][i9]), .B(multi9[24][i9]), .Out(sum9[22][i9]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum9[21][i9]), .B(sum9[22][i9]), .Out(sum9[23][i9]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum9[23][i9]), .B(feature1Bias), .Out(data_11_array[j9][i9]));
    end
  endgenerate
  
  ////ROW 10
  generate
    localparam integer j10 = 10;
    for (i10 = 0; i10 < 24; i10 = i10 + 1)
    begin: addbit10
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j10+0][i10+0]), .Out(multi10[0][i10]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j10+0][i10+1]), .Out(multi10[1][i10]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j10+0][i10+2]), .Out(multi10[2][i10]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j10+0][i10+3]), .Out(multi10[3][i10]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j10+0][i10+4]), .Out(multi10[4][i10]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j10+1][i10+0]), .Out(multi10[5][i10]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j10+1][i10+1]), .Out(multi10[6][i10]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j10+1][i10+2]), .Out(multi10[7][i10]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j10+1][i10+3]), .Out(multi10[8][i10]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j10+1][i10+4]), .Out(multi10[9][i10]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j10+2][i10+0]), .Out(multi10[10][i10]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j10+2][i10+1]), .Out(multi10[11][i10]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j10+2][i10+2]), .Out(multi10[12][i10]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j10+2][i10+3]), .Out(multi10[13][i10]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j10+2][i10+4]), .Out(multi10[14][i10]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j10+3][i10+0]), .Out(multi10[15][i10]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j10+3][i10+1]), .Out(multi10[16][i10]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j10+3][i10+2]), .Out(multi10[17][i10]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j10+3][i10+3]), .Out(multi10[18][i10]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j10+3][i10+4]), .Out(multi10[19][i10]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j10+4][i10+0]), .Out(multi10[20][i10]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j10+4][i10+1]), .Out(multi10[21][i10]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j10+4][i10+2]), .Out(multi10[22][i10]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j10+4][i10+3]), .Out(multi10[23][i10]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j10+4][i10+4]), .Out(multi10[24][i10]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi10[0][i10]), .B(multi10[1][i10]), .Out(sum10[0][i10]));
      FP16_Add stage026(.A(multi10[2][i10]), .B(multi10[3][i10]), .Out(sum10[1][i10]));
      FP16_Add stage027(.A(multi10[4][i10]), .B(multi10[5][i10]), .Out(sum10[2][i10]));
      FP16_Add stage028(.A(multi10[6][i10]), .B(multi10[7][i10]), .Out(sum10[3][i10]));
      FP16_Add stage029(.A(multi10[8][i10]), .B(multi10[9][i10]), .Out(sum10[4][i10]));
      FP16_Add stage030(.A(multi10[10][i10]), .B(multi10[11][i10]), .Out(sum10[5][i10]));
      FP16_Add stage031(.A(multi10[12][i10]), .B(multi10[13][i10]), .Out(sum10[6][i10]));
      FP16_Add stage032(.A(multi10[14][i10]), .B(multi10[15][i10]), .Out(sum10[7][i10]));
      FP16_Add stage033(.A(multi10[16][i10]), .B(multi10[17][i10]), .Out(sum10[8][i10]));
      FP16_Add stage034(.A(multi10[18][i10]), .B(multi10[19][i10]), .Out(sum10[9][i10]));
      FP16_Add stage035(.A(multi10[20][i10]), .B(multi10[21][i10]), .Out(sum10[10][i10]));
      FP16_Add stage036(.A(multi10[22][i10]), .B(multi10[23][i10]), .Out(sum10[11][i10]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum10[0][i10]), .B(sum10[1][i10]), .Out(sum10[12][i10]));
      FP16_Add stage038(.A(sum10[2][i10]), .B(sum10[3][i10]), .Out(sum10[13][i10]));
      FP16_Add stage039(.A(sum10[4][i10]), .B(sum10[5][i10]), .Out(sum10[14][i10]));
      FP16_Add stage040(.A(sum10[6][i10]), .B(sum10[7][i10]), .Out(sum10[15][i10]));
      FP16_Add stage041(.A(sum10[8][i10]), .B(sum10[9][i10]), .Out(sum10[16][i10]));
      FP16_Add stage042(.A(sum10[10][i10]), .B(sum10[11][i10]), .Out(sum10[17][i10]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum10[12][i10]), .B(sum10[13][i10]), .Out(sum10[18][i10]));
      FP16_Add stage044(.A(sum10[14][i10]), .B(sum10[15][i10]), .Out(sum10[19][i10]));
      FP16_Add stage045(.A(sum10[16][i10]), .B(sum10[17][i10]), .Out(sum10[20][i10]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum10[18][i10]), .B(sum10[19][i10]), .Out(sum10[21][i10]));
      FP16_Add stage047(.A(sum10[20][i10]), .B(multi10[24][i10]), .Out(sum10[22][i10]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum10[21][i10]), .B(sum10[22][i10]), .Out(sum10[23][i10]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum10[23][i10]), .B(feature1Bias), .Out(data_11_array[j10][i10]));
    end
  endgenerate
  
    ////ROW 11
  generate
    localparam integer j11 = 11;
    for (i11 = 0; i11 < 24; i11 = i11 + 1)
    begin: addbit11
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j11+0][i11+0]), .Out(multi11[0][i11]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j11+0][i11+1]), .Out(multi11[1][i11]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j11+0][i11+2]), .Out(multi11[2][i11]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j11+0][i11+3]), .Out(multi11[3][i11]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j11+0][i11+4]), .Out(multi11[4][i11]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j11+1][i11+0]), .Out(multi11[5][i11]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j11+1][i11+1]), .Out(multi11[6][i11]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j11+1][i11+2]), .Out(multi11[7][i11]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j11+1][i11+3]), .Out(multi11[8][i11]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j11+1][i11+4]), .Out(multi11[9][i11]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j11+2][i11+0]), .Out(multi11[10][i11]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j11+2][i11+1]), .Out(multi11[11][i11]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j11+2][i11+2]), .Out(multi11[12][i11]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j11+2][i11+3]), .Out(multi11[13][i11]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j11+2][i11+4]), .Out(multi11[14][i11]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j11+3][i11+0]), .Out(multi11[15][i11]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j11+3][i11+1]), .Out(multi11[16][i11]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j11+3][i11+2]), .Out(multi11[17][i11]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j11+3][i11+3]), .Out(multi11[18][i11]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j11+3][i11+4]), .Out(multi11[19][i11]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j11+4][i11+0]), .Out(multi11[20][i11]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j11+4][i11+1]), .Out(multi11[21][i11]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j11+4][i11+2]), .Out(multi11[22][i11]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j11+4][i11+3]), .Out(multi11[23][i11]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j11+4][i11+4]), .Out(multi11[24][i11]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi11[0][i11]), .B(multi11[1][i11]), .Out(sum11[0][i11]));
      FP16_Add stage026(.A(multi11[2][i11]), .B(multi11[3][i11]), .Out(sum11[1][i11]));
      FP16_Add stage027(.A(multi11[4][i11]), .B(multi11[5][i11]), .Out(sum11[2][i11]));
      FP16_Add stage028(.A(multi11[6][i11]), .B(multi11[7][i11]), .Out(sum11[3][i11]));
      FP16_Add stage029(.A(multi11[8][i11]), .B(multi11[9][i11]), .Out(sum11[4][i11]));
      FP16_Add stage030(.A(multi11[10][i11]), .B(multi11[11][i11]), .Out(sum11[5][i11]));
      FP16_Add stage031(.A(multi11[12][i11]), .B(multi11[13][i11]), .Out(sum11[6][i11]));
      FP16_Add stage032(.A(multi11[14][i11]), .B(multi11[15][i11]), .Out(sum11[7][i11]));
      FP16_Add stage033(.A(multi11[16][i11]), .B(multi11[17][i11]), .Out(sum11[8][i11]));
      FP16_Add stage034(.A(multi11[18][i11]), .B(multi11[19][i11]), .Out(sum11[9][i11]));
      FP16_Add stage035(.A(multi11[20][i11]), .B(multi11[21][i11]), .Out(sum11[10][i11]));
      FP16_Add stage036(.A(multi11[22][i11]), .B(multi11[23][i11]), .Out(sum11[11][i11]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum11[0][i11]), .B(sum11[1][i11]), .Out(sum11[12][i11]));
      FP16_Add stage038(.A(sum11[2][i11]), .B(sum11[3][i11]), .Out(sum11[13][i11]));
      FP16_Add stage039(.A(sum11[4][i11]), .B(sum11[5][i11]), .Out(sum11[14][i11]));
      FP16_Add stage040(.A(sum11[6][i11]), .B(sum11[7][i11]), .Out(sum11[15][i11]));
      FP16_Add stage041(.A(sum11[8][i11]), .B(sum11[9][i11]), .Out(sum11[16][i11]));
      FP16_Add stage042(.A(sum11[10][i11]), .B(sum11[11][i11]), .Out(sum11[17][i11]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum11[12][i11]), .B(sum11[13][i11]), .Out(sum11[18][i11]));
      FP16_Add stage044(.A(sum11[14][i11]), .B(sum11[15][i11]), .Out(sum11[19][i11]));
      FP16_Add stage045(.A(sum11[16][i11]), .B(sum11[17][i11]), .Out(sum11[20][i11]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum11[18][i11]), .B(sum11[19][i11]), .Out(sum11[21][i11]));
      FP16_Add stage047(.A(sum11[20][i11]), .B(multi11[24][i11]), .Out(sum11[22][i11]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum11[21][i11]), .B(sum11[22][i11]), .Out(sum11[23][i11]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum11[23][i11]), .B(feature1Bias), .Out(data_11_array[j11][i11]));
    end
  endgenerate

  ////ROW 12
  generate
    localparam integer j12 = 12;
    for (i12 = 0; i12 < 24; i12 = i12 + 1)
    begin: addbit12
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j12+0][i12+0]), .Out(multi12[0][i12]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j12+0][i12+1]), .Out(multi12[1][i12]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j12+0][i12+2]), .Out(multi12[2][i12]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j12+0][i12+3]), .Out(multi12[3][i12]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j12+0][i12+4]), .Out(multi12[4][i12]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j12+1][i12+0]), .Out(multi12[5][i12]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j12+1][i12+1]), .Out(multi12[6][i12]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j12+1][i12+2]), .Out(multi12[7][i12]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j12+1][i12+3]), .Out(multi12[8][i12]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j12+1][i12+4]), .Out(multi12[9][i12]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j12+2][i12+0]), .Out(multi12[10][i12]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j12+2][i12+1]), .Out(multi12[11][i12]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j12+2][i12+2]), .Out(multi12[12][i12]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j12+2][i12+3]), .Out(multi12[13][i12]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j12+2][i12+4]), .Out(multi12[14][i12]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j12+3][i12+0]), .Out(multi12[15][i12]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j12+3][i12+1]), .Out(multi12[16][i12]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j12+3][i12+2]), .Out(multi12[17][i12]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j12+3][i12+3]), .Out(multi12[18][i12]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j12+3][i12+4]), .Out(multi12[19][i12]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j12+4][i12+0]), .Out(multi12[20][i12]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j12+4][i12+1]), .Out(multi12[21][i12]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j12+4][i12+2]), .Out(multi12[22][i12]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j12+4][i12+3]), .Out(multi12[23][i12]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j12+4][i12+4]), .Out(multi12[24][i12]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi12[0][i12]), .B(multi12[1][i12]), .Out(sum12[0][i12]));
      FP16_Add stage026(.A(multi12[2][i12]), .B(multi12[3][i12]), .Out(sum12[1][i12]));
      FP16_Add stage027(.A(multi12[4][i12]), .B(multi12[5][i12]), .Out(sum12[2][i12]));
      FP16_Add stage028(.A(multi12[6][i12]), .B(multi12[7][i12]), .Out(sum12[3][i12]));
      FP16_Add stage029(.A(multi12[8][i12]), .B(multi12[9][i12]), .Out(sum12[4][i12]));
      FP16_Add stage030(.A(multi12[10][i12]), .B(multi12[11][i12]), .Out(sum12[5][i12]));
      FP16_Add stage031(.A(multi12[12][i12]), .B(multi12[13][i12]), .Out(sum12[6][i12]));
      FP16_Add stage032(.A(multi12[14][i12]), .B(multi12[15][i12]), .Out(sum12[7][i12]));
      FP16_Add stage033(.A(multi12[16][i12]), .B(multi12[17][i12]), .Out(sum12[8][i12]));
      FP16_Add stage034(.A(multi12[18][i12]), .B(multi12[19][i12]), .Out(sum12[9][i12]));
      FP16_Add stage035(.A(multi12[20][i12]), .B(multi12[21][i12]), .Out(sum12[10][i12]));
      FP16_Add stage036(.A(multi12[22][i12]), .B(multi12[23][i12]), .Out(sum12[11][i12]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum12[0][i12]), .B(sum12[1][i12]), .Out(sum12[12][i12]));
      FP16_Add stage038(.A(sum12[2][i12]), .B(sum12[3][i12]), .Out(sum12[13][i12]));
      FP16_Add stage039(.A(sum12[4][i12]), .B(sum12[5][i12]), .Out(sum12[14][i12]));
      FP16_Add stage040(.A(sum12[6][i12]), .B(sum12[7][i12]), .Out(sum12[15][i12]));
      FP16_Add stage041(.A(sum12[8][i12]), .B(sum12[9][i12]), .Out(sum12[16][i12]));
      FP16_Add stage042(.A(sum12[10][i12]), .B(sum12[11][i12]), .Out(sum12[17][i12]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum12[12][i12]), .B(sum12[13][i12]), .Out(sum12[18][i12]));
      FP16_Add stage044(.A(sum12[14][i12]), .B(sum12[15][i12]), .Out(sum12[19][i12]));
      FP16_Add stage045(.A(sum12[16][i12]), .B(sum12[17][i12]), .Out(sum12[20][i12]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum12[18][i12]), .B(sum12[19][i12]), .Out(sum12[21][i12]));
      FP16_Add stage047(.A(sum12[20][i12]), .B(multi12[24][i12]), .Out(sum12[22][i12]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum12[21][i12]), .B(sum12[22][i12]), .Out(sum12[23][i12]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum12[23][i12]), .B(feature1Bias), .Out(data_11_array[j12][i12]));
    end
  endgenerate

  ////ROW 13
  generate
    localparam integer j13 = 13;
    for (i13 = 0; i13 < 24; i13 = i13 + 1)
    begin: addbit13
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j13+0][i13+0]), .Out(multi13[0][i13]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j13+0][i13+1]), .Out(multi13[1][i13]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j13+0][i13+2]), .Out(multi13[2][i13]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j13+0][i13+3]), .Out(multi13[3][i13]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j13+0][i13+4]), .Out(multi13[4][i13]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j13+1][i13+0]), .Out(multi13[5][i13]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j13+1][i13+1]), .Out(multi13[6][i13]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j13+1][i13+2]), .Out(multi13[7][i13]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j13+1][i13+3]), .Out(multi13[8][i13]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j13+1][i13+4]), .Out(multi13[9][i13]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j13+2][i13+0]), .Out(multi13[10][i13]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j13+2][i13+1]), .Out(multi13[11][i13]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j13+2][i13+2]), .Out(multi13[12][i13]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j13+2][i13+3]), .Out(multi13[13][i13]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j13+2][i13+4]), .Out(multi13[14][i13]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j13+3][i13+0]), .Out(multi13[15][i13]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j13+3][i13+1]), .Out(multi13[16][i13]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j13+3][i13+2]), .Out(multi13[17][i13]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j13+3][i13+3]), .Out(multi13[18][i13]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j13+3][i13+4]), .Out(multi13[19][i13]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j13+4][i13+0]), .Out(multi13[20][i13]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j13+4][i13+1]), .Out(multi13[21][i13]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j13+4][i13+2]), .Out(multi13[22][i13]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j13+4][i13+3]), .Out(multi13[23][i13]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j13+4][i13+4]), .Out(multi13[24][i13]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi13[0][i13]), .B(multi13[1][i13]), .Out(sum13[0][i13]));
      FP16_Add stage026(.A(multi13[2][i13]), .B(multi13[3][i13]), .Out(sum13[1][i13]));
      FP16_Add stage027(.A(multi13[4][i13]), .B(multi13[5][i13]), .Out(sum13[2][i13]));
      FP16_Add stage028(.A(multi13[6][i13]), .B(multi13[7][i13]), .Out(sum13[3][i13]));
      FP16_Add stage029(.A(multi13[8][i13]), .B(multi13[9][i13]), .Out(sum13[4][i13]));
      FP16_Add stage030(.A(multi13[10][i13]), .B(multi13[11][i13]), .Out(sum13[5][i13]));
      FP16_Add stage031(.A(multi13[12][i13]), .B(multi13[13][i13]), .Out(sum13[6][i13]));
      FP16_Add stage032(.A(multi13[14][i13]), .B(multi13[15][i13]), .Out(sum13[7][i13]));
      FP16_Add stage033(.A(multi13[16][i13]), .B(multi13[17][i13]), .Out(sum13[8][i13]));
      FP16_Add stage034(.A(multi13[18][i13]), .B(multi13[19][i13]), .Out(sum13[9][i13]));
      FP16_Add stage035(.A(multi13[20][i13]), .B(multi13[21][i13]), .Out(sum13[10][i13]));
      FP16_Add stage036(.A(multi13[22][i13]), .B(multi13[23][i13]), .Out(sum13[11][i13]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum13[0][i13]), .B(sum13[1][i13]), .Out(sum13[12][i13]));
      FP16_Add stage038(.A(sum13[2][i13]), .B(sum13[3][i13]), .Out(sum13[13][i13]));
      FP16_Add stage039(.A(sum13[4][i13]), .B(sum13[5][i13]), .Out(sum13[14][i13]));
      FP16_Add stage040(.A(sum13[6][i13]), .B(sum13[7][i13]), .Out(sum13[15][i13]));
      FP16_Add stage041(.A(sum13[8][i13]), .B(sum13[9][i13]), .Out(sum13[16][i13]));
      FP16_Add stage042(.A(sum13[10][i13]), .B(sum13[11][i13]), .Out(sum13[17][i13]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum13[12][i13]), .B(sum13[13][i13]), .Out(sum13[18][i13]));
      FP16_Add stage044(.A(sum13[14][i13]), .B(sum13[15][i13]), .Out(sum13[19][i13]));
      FP16_Add stage045(.A(sum13[16][i13]), .B(sum13[17][i13]), .Out(sum13[20][i13]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum13[18][i13]), .B(sum13[19][i13]), .Out(sum13[21][i13]));
      FP16_Add stage047(.A(sum13[20][i13]), .B(multi13[24][i13]), .Out(sum13[22][i13]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum13[21][i13]), .B(sum13[22][i13]), .Out(sum13[23][i13]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum13[23][i13]), .B(feature1Bias), .Out(data_11_array[j13][i13]));
    end
  endgenerate

  ////ROW 014
  generate
    localparam integer j14 = 14;
    for (i14 = 0; i14 < 24; i14 = i14 + 1)
    begin: addbit14
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j14+0][i14+0]), .Out(multi14[0][i14]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j14+0][i14+1]), .Out(multi14[1][i14]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j14+0][i14+2]), .Out(multi14[2][i14]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j14+0][i14+3]), .Out(multi14[3][i14]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j14+0][i14+4]), .Out(multi14[4][i14]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j14+1][i14+0]), .Out(multi14[5][i14]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j14+1][i14+1]), .Out(multi14[6][i14]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j14+1][i14+2]), .Out(multi14[7][i14]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j14+1][i14+3]), .Out(multi14[8][i14]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j14+1][i14+4]), .Out(multi14[9][i14]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j14+2][i14+0]), .Out(multi14[10][i14]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j14+2][i14+1]), .Out(multi14[11][i14]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j14+2][i14+2]), .Out(multi14[12][i14]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j14+2][i14+3]), .Out(multi14[13][i14]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j14+2][i14+4]), .Out(multi14[14][i14]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j14+3][i14+0]), .Out(multi14[15][i14]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j14+3][i14+1]), .Out(multi14[16][i14]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j14+3][i14+2]), .Out(multi14[17][i14]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j14+3][i14+3]), .Out(multi14[18][i14]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j14+3][i14+4]), .Out(multi14[19][i14]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j14+4][i14+0]), .Out(multi14[20][i14]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j14+4][i14+1]), .Out(multi14[21][i14]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j14+4][i14+2]), .Out(multi14[22][i14]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j14+4][i14+3]), .Out(multi14[23][i14]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j14+4][i14+4]), .Out(multi14[24][i14]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi14[0][i14]), .B(multi14[1][i14]), .Out(sum14[0][i14]));
      FP16_Add stage026(.A(multi14[2][i14]), .B(multi14[3][i14]), .Out(sum14[1][i14]));
      FP16_Add stage027(.A(multi14[4][i14]), .B(multi14[5][i14]), .Out(sum14[2][i14]));
      FP16_Add stage028(.A(multi14[6][i14]), .B(multi14[7][i14]), .Out(sum14[3][i14]));
      FP16_Add stage029(.A(multi14[8][i14]), .B(multi14[9][i14]), .Out(sum14[4][i14]));
      FP16_Add stage030(.A(multi14[10][i14]), .B(multi14[11][i14]), .Out(sum14[5][i14]));
      FP16_Add stage031(.A(multi14[12][i14]), .B(multi14[13][i14]), .Out(sum14[6][i14]));
      FP16_Add stage032(.A(multi14[14][i14]), .B(multi14[15][i14]), .Out(sum14[7][i14]));
      FP16_Add stage033(.A(multi14[16][i14]), .B(multi14[17][i14]), .Out(sum14[8][i14]));
      FP16_Add stage034(.A(multi14[18][i14]), .B(multi14[19][i14]), .Out(sum14[9][i14]));
      FP16_Add stage035(.A(multi14[20][i14]), .B(multi14[21][i14]), .Out(sum14[10][i14]));
      FP16_Add stage036(.A(multi14[22][i14]), .B(multi14[23][i14]), .Out(sum14[11][i14]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum14[0][i14]), .B(sum14[1][i14]), .Out(sum14[12][i14]));
      FP16_Add stage038(.A(sum14[2][i14]), .B(sum14[3][i14]), .Out(sum14[13][i14]));
      FP16_Add stage039(.A(sum14[4][i14]), .B(sum14[5][i14]), .Out(sum14[14][i14]));
      FP16_Add stage040(.A(sum14[6][i14]), .B(sum14[7][i14]), .Out(sum14[15][i14]));
      FP16_Add stage041(.A(sum14[8][i14]), .B(sum14[9][i14]), .Out(sum14[16][i14]));
      FP16_Add stage042(.A(sum14[10][i14]), .B(sum14[11][i14]), .Out(sum14[17][i14]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum14[12][i14]), .B(sum14[13][i14]), .Out(sum14[18][i14]));
      FP16_Add stage044(.A(sum14[14][i14]), .B(sum14[15][i14]), .Out(sum14[19][i14]));
      FP16_Add stage045(.A(sum14[16][i14]), .B(sum14[17][i14]), .Out(sum14[20][i14]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum14[18][i14]), .B(sum14[19][i14]), .Out(sum14[21][i14]));
      FP16_Add stage047(.A(sum14[20][i14]), .B(multi14[24][i14]), .Out(sum14[22][i14]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum14[21][i14]), .B(sum14[22][i14]), .Out(sum14[23][i14]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum14[23][i14]), .B(feature1Bias), .Out(data_11_array[j14][i14]));
    end
  endgenerate

  ////ROW 15
  generate
    localparam integer j15 = 15;
    for (i15 = 0; i15 < 24; i15 = i15 + 1)
    begin: addbit15
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j15+0][i15+0]), .Out(multi15[0][i15]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j15+0][i15+1]), .Out(multi15[1][i15]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j15+0][i15+2]), .Out(multi15[2][i15]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j15+0][i15+3]), .Out(multi15[3][i15]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j15+0][i15+4]), .Out(multi15[4][i15]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j15+1][i15+0]), .Out(multi15[5][i15]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j15+1][i15+1]), .Out(multi15[6][i15]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j15+1][i15+2]), .Out(multi15[7][i15]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j15+1][i15+3]), .Out(multi15[8][i15]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j15+1][i15+4]), .Out(multi15[9][i15]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j15+2][i15+0]), .Out(multi15[10][i15]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j15+2][i15+1]), .Out(multi15[11][i15]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j15+2][i15+2]), .Out(multi15[12][i15]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j15+2][i15+3]), .Out(multi15[13][i15]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j15+2][i15+4]), .Out(multi15[14][i15]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j15+3][i15+0]), .Out(multi15[15][i15]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j15+3][i15+1]), .Out(multi15[16][i15]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j15+3][i15+2]), .Out(multi15[17][i15]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j15+3][i15+3]), .Out(multi15[18][i15]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j15+3][i15+4]), .Out(multi15[19][i15]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j15+4][i15+0]), .Out(multi15[20][i15]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j15+4][i15+1]), .Out(multi15[21][i15]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j15+4][i15+2]), .Out(multi15[22][i15]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j15+4][i15+3]), .Out(multi15[23][i15]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j15+4][i15+4]), .Out(multi15[24][i15]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi15[0][i15]), .B(multi15[1][i15]), .Out(sum15[0][i15]));
      FP16_Add stage026(.A(multi15[2][i15]), .B(multi15[3][i15]), .Out(sum15[1][i15]));
      FP16_Add stage027(.A(multi15[4][i15]), .B(multi15[5][i15]), .Out(sum15[2][i15]));
      FP16_Add stage028(.A(multi15[6][i15]), .B(multi15[7][i15]), .Out(sum15[3][i15]));
      FP16_Add stage029(.A(multi15[8][i15]), .B(multi15[9][i15]), .Out(sum15[4][i15]));
      FP16_Add stage030(.A(multi15[10][i15]), .B(multi15[11][i15]), .Out(sum15[5][i15]));
      FP16_Add stage031(.A(multi15[12][i15]), .B(multi15[13][i15]), .Out(sum15[6][i15]));
      FP16_Add stage032(.A(multi15[14][i15]), .B(multi15[15][i15]), .Out(sum15[7][i15]));
      FP16_Add stage033(.A(multi15[16][i15]), .B(multi15[17][i15]), .Out(sum15[8][i15]));
      FP16_Add stage034(.A(multi15[18][i15]), .B(multi15[19][i15]), .Out(sum15[9][i15]));
      FP16_Add stage035(.A(multi15[20][i15]), .B(multi15[21][i15]), .Out(sum15[10][i15]));
      FP16_Add stage036(.A(multi15[22][i15]), .B(multi15[23][i15]), .Out(sum15[11][i15]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum15[0][i15]), .B(sum15[1][i15]), .Out(sum15[12][i15]));
      FP16_Add stage038(.A(sum15[2][i15]), .B(sum15[3][i15]), .Out(sum15[13][i15]));
      FP16_Add stage039(.A(sum15[4][i15]), .B(sum15[5][i15]), .Out(sum15[14][i15]));
      FP16_Add stage040(.A(sum15[6][i15]), .B(sum15[7][i15]), .Out(sum15[15][i15]));
      FP16_Add stage041(.A(sum15[8][i15]), .B(sum15[9][i15]), .Out(sum15[16][i15]));
      FP16_Add stage042(.A(sum15[10][i15]), .B(sum15[11][i15]), .Out(sum15[17][i15]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum15[12][i15]), .B(sum15[13][i15]), .Out(sum15[18][i15]));
      FP16_Add stage044(.A(sum15[14][i15]), .B(sum15[15][i15]), .Out(sum15[19][i15]));
      FP16_Add stage045(.A(sum15[16][i15]), .B(sum15[17][i15]), .Out(sum15[20][i15]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum15[18][i15]), .B(sum15[19][i15]), .Out(sum15[21][i15]));
      FP16_Add stage047(.A(sum15[20][i15]), .B(multi15[24][i15]), .Out(sum15[22][i15]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum15[21][i15]), .B(sum15[22][i15]), .Out(sum15[23][i15]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum15[23][i15]), .B(feature1Bias), .Out(data_11_array[j15][i15]));
    end
  endgenerate
  
  ////ROW 16
  generate
    localparam integer j16 = 16;
    for (i16 = 0; i16 < 24; i16 = i16 + 1)
    begin: addbit16
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j16+0][i16+0]), .Out(multi16[0][i16]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j16+0][i16+1]), .Out(multi16[1][i16]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j16+0][i16+2]), .Out(multi16[2][i16]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j16+0][i16+3]), .Out(multi16[3][i16]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j16+0][i16+4]), .Out(multi16[4][i16]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j16+1][i16+0]), .Out(multi16[5][i16]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j16+1][i16+1]), .Out(multi16[6][i16]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j16+1][i16+2]), .Out(multi16[7][i16]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j16+1][i16+3]), .Out(multi16[8][i16]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j16+1][i16+4]), .Out(multi16[9][i16]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j16+2][i16+0]), .Out(multi16[10][i16]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j16+2][i16+1]), .Out(multi16[11][i16]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j16+2][i16+2]), .Out(multi16[12][i16]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j16+2][i16+3]), .Out(multi16[13][i16]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j16+2][i16+4]), .Out(multi16[14][i16]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j16+3][i16+0]), .Out(multi16[15][i16]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j16+3][i16+1]), .Out(multi16[16][i16]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j16+3][i16+2]), .Out(multi16[17][i16]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j16+3][i16+3]), .Out(multi16[18][i16]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j16+3][i16+4]), .Out(multi16[19][i16]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j16+4][i16+0]), .Out(multi16[20][i16]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j16+4][i16+1]), .Out(multi16[21][i16]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j16+4][i16+2]), .Out(multi16[22][i16]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j16+4][i16+3]), .Out(multi16[23][i16]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j16+4][i16+4]), .Out(multi16[24][i16]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi16[0][i16]), .B(multi16[1][i16]), .Out(sum16[0][i16]));
      FP16_Add stage026(.A(multi16[2][i16]), .B(multi16[3][i16]), .Out(sum16[1][i16]));
      FP16_Add stage027(.A(multi16[4][i16]), .B(multi16[5][i16]), .Out(sum16[2][i16]));
      FP16_Add stage028(.A(multi16[6][i16]), .B(multi16[7][i16]), .Out(sum16[3][i16]));
      FP16_Add stage029(.A(multi16[8][i16]), .B(multi16[9][i16]), .Out(sum16[4][i16]));
      FP16_Add stage030(.A(multi16[10][i16]), .B(multi16[11][i16]), .Out(sum16[5][i16]));
      FP16_Add stage031(.A(multi16[12][i16]), .B(multi16[13][i16]), .Out(sum16[6][i16]));
      FP16_Add stage032(.A(multi16[14][i16]), .B(multi16[15][i16]), .Out(sum16[7][i16]));
      FP16_Add stage033(.A(multi16[16][i16]), .B(multi16[17][i16]), .Out(sum16[8][i16]));
      FP16_Add stage034(.A(multi16[18][i16]), .B(multi16[19][i16]), .Out(sum16[9][i16]));
      FP16_Add stage035(.A(multi16[20][i16]), .B(multi16[21][i16]), .Out(sum16[10][i16]));
      FP16_Add stage036(.A(multi16[22][i16]), .B(multi16[23][i16]), .Out(sum16[11][i16]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum16[0][i16]), .B(sum16[1][i16]), .Out(sum16[12][i16]));
      FP16_Add stage038(.A(sum16[2][i16]), .B(sum16[3][i16]), .Out(sum16[13][i16]));
      FP16_Add stage039(.A(sum16[4][i16]), .B(sum16[5][i16]), .Out(sum16[14][i16]));
      FP16_Add stage040(.A(sum16[6][i16]), .B(sum16[7][i16]), .Out(sum16[15][i16]));
      FP16_Add stage041(.A(sum16[8][i16]), .B(sum16[9][i16]), .Out(sum16[16][i16]));
      FP16_Add stage042(.A(sum16[10][i16]), .B(sum16[11][i16]), .Out(sum16[17][i16]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum16[12][i16]), .B(sum16[13][i16]), .Out(sum16[18][i16]));
      FP16_Add stage044(.A(sum16[14][i16]), .B(sum16[15][i16]), .Out(sum16[19][i16]));
      FP16_Add stage045(.A(sum16[16][i16]), .B(sum16[17][i16]), .Out(sum16[20][i16]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum16[18][i16]), .B(sum16[19][i16]), .Out(sum16[21][i16]));
      FP16_Add stage047(.A(sum16[20][i16]), .B(multi16[24][i16]), .Out(sum16[22][i16]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum16[21][i16]), .B(sum16[22][i16]), .Out(sum16[23][i16]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum16[23][i16]), .B(feature1Bias), .Out(data_11_array[j16][i16]));
    end
  endgenerate
  
  ////ROW 17
  generate
    localparam integer j17 = 17;
    for (i17 = 0; i17 < 24; i17 = i17 + 1)
    begin: addbit17
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j17+0][i17+0]), .Out(multi17[0][i17]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j17+0][i17+1]), .Out(multi17[1][i17]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j17+0][i17+2]), .Out(multi17[2][i17]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j17+0][i17+3]), .Out(multi17[3][i17]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j17+0][i17+4]), .Out(multi17[4][i17]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j17+1][i17+0]), .Out(multi17[5][i17]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j17+1][i17+1]), .Out(multi17[6][i17]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j17+1][i17+2]), .Out(multi17[7][i17]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j17+1][i17+3]), .Out(multi17[8][i17]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j17+1][i17+4]), .Out(multi17[9][i17]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j17+2][i17+0]), .Out(multi17[10][i17]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j17+2][i17+1]), .Out(multi17[11][i17]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j17+2][i17+2]), .Out(multi17[12][i17]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j17+2][i17+3]), .Out(multi17[13][i17]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j17+2][i17+4]), .Out(multi17[14][i17]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j17+3][i17+0]), .Out(multi17[15][i17]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j17+3][i17+1]), .Out(multi17[16][i17]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j17+3][i17+2]), .Out(multi17[17][i17]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j17+3][i17+3]), .Out(multi17[18][i17]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j17+3][i17+4]), .Out(multi17[19][i17]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j17+4][i17+0]), .Out(multi17[20][i17]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j17+4][i17+1]), .Out(multi17[21][i17]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j17+4][i17+2]), .Out(multi17[22][i17]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j17+4][i17+3]), .Out(multi17[23][i17]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j17+4][i17+4]), .Out(multi17[24][i17]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi17[0][i17]), .B(multi17[1][i17]), .Out(sum17[0][i17]));
      FP16_Add stage026(.A(multi17[2][i17]), .B(multi17[3][i17]), .Out(sum17[1][i17]));
      FP16_Add stage027(.A(multi17[4][i17]), .B(multi17[5][i17]), .Out(sum17[2][i17]));
      FP16_Add stage028(.A(multi17[6][i17]), .B(multi17[7][i17]), .Out(sum17[3][i17]));
      FP16_Add stage029(.A(multi17[8][i17]), .B(multi17[9][i17]), .Out(sum17[4][i17]));
      FP16_Add stage030(.A(multi17[10][i17]), .B(multi17[11][i17]), .Out(sum17[5][i17]));
      FP16_Add stage031(.A(multi17[12][i17]), .B(multi17[13][i17]), .Out(sum17[6][i17]));
      FP16_Add stage032(.A(multi17[14][i17]), .B(multi17[15][i17]), .Out(sum17[7][i17]));
      FP16_Add stage033(.A(multi17[16][i17]), .B(multi17[17][i17]), .Out(sum17[8][i17]));
      FP16_Add stage034(.A(multi17[18][i17]), .B(multi17[19][i17]), .Out(sum17[9][i17]));
      FP16_Add stage035(.A(multi17[20][i17]), .B(multi17[21][i17]), .Out(sum17[10][i17]));
      FP16_Add stage036(.A(multi17[22][i17]), .B(multi17[23][i17]), .Out(sum17[11][i17]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum17[0][i17]), .B(sum17[1][i17]), .Out(sum17[12][i17]));
      FP16_Add stage038(.A(sum17[2][i17]), .B(sum17[3][i17]), .Out(sum17[13][i17]));
      FP16_Add stage039(.A(sum17[4][i17]), .B(sum17[5][i17]), .Out(sum17[14][i17]));
      FP16_Add stage040(.A(sum17[6][i17]), .B(sum17[7][i17]), .Out(sum17[15][i17]));
      FP16_Add stage041(.A(sum17[8][i17]), .B(sum17[9][i17]), .Out(sum17[16][i17]));
      FP16_Add stage042(.A(sum17[10][i17]), .B(sum17[11][i17]), .Out(sum17[17][i17]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum17[12][i17]), .B(sum17[13][i17]), .Out(sum17[18][i17]));
      FP16_Add stage044(.A(sum17[14][i17]), .B(sum17[15][i17]), .Out(sum17[19][i17]));
      FP16_Add stage045(.A(sum17[16][i17]), .B(sum17[17][i17]), .Out(sum17[20][i17]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum17[18][i17]), .B(sum17[19][i17]), .Out(sum17[21][i17]));
      FP16_Add stage047(.A(sum17[20][i17]), .B(multi17[24][i17]), .Out(sum17[22][i17]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum17[21][i17]), .B(sum17[22][i17]), .Out(sum17[23][i17]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum17[23][i17]), .B(feature1Bias), .Out(data_11_array[j17][i17]));
    end
  endgenerate

////ROW 18
  generate
    localparam integer j18 = 18;
    for (i18 = 0; i18 < 24; i18 = i18 + 1)
    begin: addbit18
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j18+0][i18+0]), .Out(multi18[0][i18]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j18+0][i18+1]), .Out(multi18[1][i18]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j18+0][i18+2]), .Out(multi18[2][i18]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j18+0][i18+3]), .Out(multi18[3][i18]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j18+0][i18+4]), .Out(multi18[4][i18]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j18+1][i18+0]), .Out(multi18[5][i18]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j18+1][i18+1]), .Out(multi18[6][i18]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j18+1][i18+2]), .Out(multi18[7][i18]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j18+1][i18+3]), .Out(multi18[8][i18]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j18+1][i18+4]), .Out(multi18[9][i18]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j18+2][i18+0]), .Out(multi18[10][i18]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j18+2][i18+1]), .Out(multi18[11][i18]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j18+2][i18+2]), .Out(multi18[12][i18]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j18+2][i18+3]), .Out(multi18[13][i18]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j18+2][i18+4]), .Out(multi18[14][i18]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j18+3][i18+0]), .Out(multi18[15][i18]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j18+3][i18+1]), .Out(multi18[16][i18]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j18+3][i18+2]), .Out(multi18[17][i18]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j18+3][i18+3]), .Out(multi18[18][i18]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j18+3][i18+4]), .Out(multi18[19][i18]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j18+4][i18+0]), .Out(multi18[20][i18]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j18+4][i18+1]), .Out(multi18[21][i18]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j18+4][i18+2]), .Out(multi18[22][i18]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j18+4][i18+3]), .Out(multi18[23][i18]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j18+4][i18+4]), .Out(multi18[24][i18]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi18[0][i18]), .B(multi18[1][i18]), .Out(sum18[0][i18]));
      FP16_Add stage026(.A(multi18[2][i18]), .B(multi18[3][i18]), .Out(sum18[1][i18]));
      FP16_Add stage027(.A(multi18[4][i18]), .B(multi18[5][i18]), .Out(sum18[2][i18]));
      FP16_Add stage028(.A(multi18[6][i18]), .B(multi18[7][i18]), .Out(sum18[3][i18]));
      FP16_Add stage029(.A(multi18[8][i18]), .B(multi18[9][i18]), .Out(sum18[4][i18]));
      FP16_Add stage030(.A(multi18[10][i18]), .B(multi18[11][i18]), .Out(sum18[5][i18]));
      FP16_Add stage031(.A(multi18[12][i18]), .B(multi18[13][i18]), .Out(sum18[6][i18]));
      FP16_Add stage032(.A(multi18[14][i18]), .B(multi18[15][i18]), .Out(sum18[7][i18]));
      FP16_Add stage033(.A(multi18[16][i18]), .B(multi18[17][i18]), .Out(sum18[8][i18]));
      FP16_Add stage034(.A(multi18[18][i18]), .B(multi18[19][i18]), .Out(sum18[9][i18]));
      FP16_Add stage035(.A(multi18[20][i18]), .B(multi18[21][i18]), .Out(sum18[10][i18]));
      FP16_Add stage036(.A(multi18[22][i18]), .B(multi18[23][i18]), .Out(sum18[11][i18]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum18[0][i18]), .B(sum18[1][i18]), .Out(sum18[12][i18]));
      FP16_Add stage038(.A(sum18[2][i18]), .B(sum18[3][i18]), .Out(sum18[13][i18]));
      FP16_Add stage039(.A(sum18[4][i18]), .B(sum18[5][i18]), .Out(sum18[14][i18]));
      FP16_Add stage040(.A(sum18[6][i18]), .B(sum18[7][i18]), .Out(sum18[15][i18]));
      FP16_Add stage041(.A(sum18[8][i18]), .B(sum18[9][i18]), .Out(sum18[16][i18]));
      FP16_Add stage042(.A(sum18[10][i18]), .B(sum18[11][i18]), .Out(sum18[17][i18]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum18[12][i18]), .B(sum18[13][i18]), .Out(sum18[18][i18]));
      FP16_Add stage044(.A(sum18[14][i18]), .B(sum18[15][i18]), .Out(sum18[19][i18]));
      FP16_Add stage045(.A(sum18[16][i18]), .B(sum18[17][i18]), .Out(sum18[20][i18]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum18[18][i18]), .B(sum18[19][i18]), .Out(sum18[21][i18]));
      FP16_Add stage047(.A(sum18[20][i18]), .B(multi18[24][i18]), .Out(sum18[22][i18]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum18[21][i18]), .B(sum18[22][i18]), .Out(sum18[23][i18]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum18[23][i18]), .B(feature1Bias), .Out(data_11_array[j18][i18]));
    end
  endgenerate

////ROW 19
  generate
    localparam integer j19 = 19;
    for (i19 = 0; i19 < 24; i19 = i19 + 1)
    begin: addbit19
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j19+0][i19+0]), .Out(multi19[0][i19]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j19+0][i19+1]), .Out(multi19[1][i19]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j19+0][i19+2]), .Out(multi19[2][i19]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j19+0][i19+3]), .Out(multi19[3][i19]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j19+0][i19+4]), .Out(multi19[4][i19]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j19+1][i19+0]), .Out(multi19[5][i19]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j19+1][i19+1]), .Out(multi19[6][i19]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j19+1][i19+2]), .Out(multi19[7][i19]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j19+1][i19+3]), .Out(multi19[8][i19]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j19+1][i19+4]), .Out(multi19[9][i19]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j19+2][i19+0]), .Out(multi19[10][i19]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j19+2][i19+1]), .Out(multi19[11][i19]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j19+2][i19+2]), .Out(multi19[12][i19]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j19+2][i19+3]), .Out(multi19[13][i19]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j19+2][i19+4]), .Out(multi19[14][i19]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j19+3][i19+0]), .Out(multi19[15][i19]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j19+3][i19+1]), .Out(multi19[16][i19]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j19+3][i19+2]), .Out(multi19[17][i19]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j19+3][i19+3]), .Out(multi19[18][i19]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j19+3][i19+4]), .Out(multi19[19][i19]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j19+4][i19+0]), .Out(multi19[20][i19]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j19+4][i19+1]), .Out(multi19[21][i19]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j19+4][i19+2]), .Out(multi19[22][i19]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j19+4][i19+3]), .Out(multi19[23][i19]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j19+4][i19+4]), .Out(multi19[24][i19]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi19[0][i19]), .B(multi19[1][i19]), .Out(sum19[0][i19]));
      FP16_Add stage026(.A(multi19[2][i19]), .B(multi19[3][i19]), .Out(sum19[1][i19]));
      FP16_Add stage027(.A(multi19[4][i19]), .B(multi19[5][i19]), .Out(sum19[2][i19]));
      FP16_Add stage028(.A(multi19[6][i19]), .B(multi19[7][i19]), .Out(sum19[3][i19]));
      FP16_Add stage029(.A(multi19[8][i19]), .B(multi19[9][i19]), .Out(sum19[4][i19]));
      FP16_Add stage030(.A(multi19[10][i19]), .B(multi19[11][i19]), .Out(sum19[5][i19]));
      FP16_Add stage031(.A(multi19[12][i19]), .B(multi19[13][i19]), .Out(sum19[6][i19]));
      FP16_Add stage032(.A(multi19[14][i19]), .B(multi19[15][i19]), .Out(sum19[7][i19]));
      FP16_Add stage033(.A(multi19[16][i19]), .B(multi19[17][i19]), .Out(sum19[8][i19]));
      FP16_Add stage034(.A(multi19[18][i19]), .B(multi19[19][i19]), .Out(sum19[9][i19]));
      FP16_Add stage035(.A(multi19[20][i19]), .B(multi19[21][i19]), .Out(sum19[10][i19]));
      FP16_Add stage036(.A(multi19[22][i19]), .B(multi19[23][i19]), .Out(sum19[11][i19]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum19[0][i19]), .B(sum19[1][i19]), .Out(sum19[12][i19]));
      FP16_Add stage038(.A(sum19[2][i19]), .B(sum19[3][i19]), .Out(sum19[13][i19]));
      FP16_Add stage039(.A(sum19[4][i19]), .B(sum19[5][i19]), .Out(sum19[14][i19]));
      FP16_Add stage040(.A(sum19[6][i19]), .B(sum19[7][i19]), .Out(sum19[15][i19]));
      FP16_Add stage041(.A(sum19[8][i19]), .B(sum19[9][i19]), .Out(sum19[16][i19]));
      FP16_Add stage042(.A(sum19[10][i19]), .B(sum19[11][i19]), .Out(sum19[17][i19]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum19[12][i19]), .B(sum19[13][i19]), .Out(sum19[18][i19]));
      FP16_Add stage044(.A(sum19[14][i19]), .B(sum19[15][i19]), .Out(sum19[19][i19]));
      FP16_Add stage045(.A(sum19[16][i19]), .B(sum19[17][i19]), .Out(sum19[20][i19]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum19[18][i19]), .B(sum19[19][i19]), .Out(sum19[21][i19]));
      FP16_Add stage047(.A(sum19[20][i19]), .B(multi19[24][i19]), .Out(sum19[22][i19]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum19[21][i19]), .B(sum19[22][i19]), .Out(sum19[23][i19]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum19[23][i19]), .B(feature1Bias), .Out(data_11_array[j19][i19]));
    end
  endgenerate

////ROW 20
  generate
    localparam integer j20 = 20;
    for (i20 = 0; i20 < 24; i20 = i20 + 1)
    begin: addbit20
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j20+0][i20+0]), .Out(multi20[0][i20]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j20+0][i20+1]), .Out(multi20[1][i20]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j20+0][i20+2]), .Out(multi20[2][i20]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j20+0][i20+3]), .Out(multi20[3][i20]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j20+0][i20+4]), .Out(multi20[4][i20]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j20+1][i20+0]), .Out(multi20[5][i20]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j20+1][i20+1]), .Out(multi20[6][i20]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j20+1][i20+2]), .Out(multi20[7][i20]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j20+1][i20+3]), .Out(multi20[8][i20]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j20+1][i20+4]), .Out(multi20[9][i20]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j20+2][i20+0]), .Out(multi20[10][i20]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j20+2][i20+1]), .Out(multi20[11][i20]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j20+2][i20+2]), .Out(multi20[12][i20]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j20+2][i20+3]), .Out(multi20[13][i20]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j20+2][i20+4]), .Out(multi20[14][i20]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j20+3][i20+0]), .Out(multi20[15][i20]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j20+3][i20+1]), .Out(multi20[16][i20]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j20+3][i20+2]), .Out(multi20[17][i20]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j20+3][i20+3]), .Out(multi20[18][i20]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j20+3][i20+4]), .Out(multi20[19][i20]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j20+4][i20+0]), .Out(multi20[20][i20]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j20+4][i20+1]), .Out(multi20[21][i20]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j20+4][i20+2]), .Out(multi20[22][i20]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j20+4][i20+3]), .Out(multi20[23][i20]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j20+4][i20+4]), .Out(multi20[24][i20]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi20[0][i20]), .B(multi20[1][i20]), .Out(sum20[0][i20]));
      FP16_Add stage026(.A(multi20[2][i20]), .B(multi20[3][i20]), .Out(sum20[1][i20]));
      FP16_Add stage027(.A(multi20[4][i20]), .B(multi20[5][i20]), .Out(sum20[2][i20]));
      FP16_Add stage028(.A(multi20[6][i20]), .B(multi20[7][i20]), .Out(sum20[3][i20]));
      FP16_Add stage029(.A(multi20[8][i20]), .B(multi20[9][i20]), .Out(sum20[4][i20]));
      FP16_Add stage030(.A(multi20[10][i20]), .B(multi20[11][i20]), .Out(sum20[5][i20]));
      FP16_Add stage031(.A(multi20[12][i20]), .B(multi20[13][i20]), .Out(sum20[6][i20]));
      FP16_Add stage032(.A(multi20[14][i20]), .B(multi20[15][i20]), .Out(sum20[7][i20]));
      FP16_Add stage033(.A(multi20[16][i20]), .B(multi20[17][i20]), .Out(sum20[8][i20]));
      FP16_Add stage034(.A(multi20[18][i20]), .B(multi20[19][i20]), .Out(sum20[9][i20]));
      FP16_Add stage035(.A(multi20[20][i20]), .B(multi20[21][i20]), .Out(sum20[10][i20]));
      FP16_Add stage036(.A(multi20[22][i20]), .B(multi20[23][i20]), .Out(sum20[11][i20]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum20[0][i20]), .B(sum20[1][i20]), .Out(sum20[12][i20]));
      FP16_Add stage038(.A(sum20[2][i20]), .B(sum20[3][i20]), .Out(sum20[13][i20]));
      FP16_Add stage039(.A(sum20[4][i20]), .B(sum20[5][i20]), .Out(sum20[14][i20]));
      FP16_Add stage040(.A(sum20[6][i20]), .B(sum20[7][i20]), .Out(sum20[15][i20]));
      FP16_Add stage041(.A(sum20[8][i20]), .B(sum20[9][i20]), .Out(sum20[16][i20]));
      FP16_Add stage042(.A(sum20[10][i20]), .B(sum20[11][i20]), .Out(sum20[17][i20]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum20[12][i20]), .B(sum20[13][i20]), .Out(sum20[18][i20]));
      FP16_Add stage044(.A(sum20[14][i20]), .B(sum20[15][i20]), .Out(sum20[19][i20]));
      FP16_Add stage045(.A(sum20[16][i20]), .B(sum20[17][i20]), .Out(sum20[20][i20]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum20[18][i20]), .B(sum20[19][i20]), .Out(sum20[21][i20]));
      FP16_Add stage047(.A(sum20[20][i20]), .B(multi20[24][i20]), .Out(sum20[22][i20]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum20[21][i20]), .B(sum20[22][i20]), .Out(sum20[23][i20]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum20[23][i20]), .B(feature1Bias), .Out(data_11_array[j20][i20]));
    end
  endgenerate

////ROW 21
  generate
    localparam integer j21 = 21;
    for (i21 = 0; i21 < 24; i21 = i21 + 1)
    begin: addbit21
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j21+0][i21+0]), .Out(multi21[0][i21]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j21+0][i21+1]), .Out(multi21[1][i21]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j21+0][i21+2]), .Out(multi21[2][i21]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j21+0][i21+3]), .Out(multi21[3][i21]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j21+0][i21+4]), .Out(multi21[4][i21]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j21+1][i21+0]), .Out(multi21[5][i21]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j21+1][i21+1]), .Out(multi21[6][i21]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j21+1][i21+2]), .Out(multi21[7][i21]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j21+1][i21+3]), .Out(multi21[8][i21]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j21+1][i21+4]), .Out(multi21[9][i21]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j21+2][i21+0]), .Out(multi21[10][i21]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j21+2][i21+1]), .Out(multi21[11][i21]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j21+2][i21+2]), .Out(multi21[12][i21]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j21+2][i21+3]), .Out(multi21[13][i21]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j21+2][i21+4]), .Out(multi21[14][i21]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j21+3][i21+0]), .Out(multi21[15][i21]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j21+3][i21+1]), .Out(multi21[16][i21]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j21+3][i21+2]), .Out(multi21[17][i21]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j21+3][i21+3]), .Out(multi21[18][i21]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j21+3][i21+4]), .Out(multi21[19][i21]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j21+4][i21+0]), .Out(multi21[20][i21]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j21+4][i21+1]), .Out(multi21[21][i21]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j21+4][i21+2]), .Out(multi21[22][i21]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j21+4][i21+3]), .Out(multi21[23][i21]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j21+4][i21+4]), .Out(multi21[24][i21]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi21[0][i21]), .B(multi21[1][i21]), .Out(sum21[0][i21]));
      FP16_Add stage026(.A(multi21[2][i21]), .B(multi21[3][i21]), .Out(sum21[1][i21]));
      FP16_Add stage027(.A(multi21[4][i21]), .B(multi21[5][i21]), .Out(sum21[2][i21]));
      FP16_Add stage028(.A(multi21[6][i21]), .B(multi21[7][i21]), .Out(sum21[3][i21]));
      FP16_Add stage029(.A(multi21[8][i21]), .B(multi21[9][i21]), .Out(sum21[4][i21]));
      FP16_Add stage030(.A(multi21[10][i21]), .B(multi21[11][i21]), .Out(sum21[5][i21]));
      FP16_Add stage031(.A(multi21[12][i21]), .B(multi21[13][i21]), .Out(sum21[6][i21]));
      FP16_Add stage032(.A(multi21[14][i21]), .B(multi21[15][i21]), .Out(sum21[7][i21]));
      FP16_Add stage033(.A(multi21[16][i21]), .B(multi21[17][i21]), .Out(sum21[8][i21]));
      FP16_Add stage034(.A(multi21[18][i21]), .B(multi21[19][i21]), .Out(sum21[9][i21]));
      FP16_Add stage035(.A(multi21[20][i21]), .B(multi21[21][i21]), .Out(sum21[10][i21]));
      FP16_Add stage036(.A(multi21[22][i21]), .B(multi21[23][i21]), .Out(sum21[11][i21]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum21[0][i21]), .B(sum21[1][i21]), .Out(sum21[12][i21]));
      FP16_Add stage038(.A(sum21[2][i21]), .B(sum21[3][i21]), .Out(sum21[13][i21]));
      FP16_Add stage039(.A(sum21[4][i21]), .B(sum21[5][i21]), .Out(sum21[14][i21]));
      FP16_Add stage040(.A(sum21[6][i21]), .B(sum21[7][i21]), .Out(sum21[15][i21]));
      FP16_Add stage041(.A(sum21[8][i21]), .B(sum21[9][i21]), .Out(sum21[16][i21]));
      FP16_Add stage042(.A(sum21[10][i21]), .B(sum21[11][i21]), .Out(sum21[17][i21]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum21[12][i21]), .B(sum21[13][i21]), .Out(sum21[18][i21]));
      FP16_Add stage044(.A(sum21[14][i21]), .B(sum21[15][i21]), .Out(sum21[19][i21]));
      FP16_Add stage045(.A(sum21[16][i21]), .B(sum21[17][i21]), .Out(sum21[20][i21]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum21[18][i21]), .B(sum21[19][i21]), .Out(sum21[21][i21]));
      FP16_Add stage047(.A(sum21[20][i21]), .B(multi21[24][i21]), .Out(sum21[22][i21]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum21[21][i21]), .B(sum21[22][i21]), .Out(sum21[23][i21]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum21[23][i21]), .B(feature1Bias), .Out(data_11_array[j21][i21]));
    end
  endgenerate

////ROW 22
  generate
    localparam integer j22 = 22;
    for (i22 = 0; i22 < 24; i22 = i22 + 1)
    begin: addbit22
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j22+0][i22+0]), .Out(multi22[0][i22]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j22+0][i22+1]), .Out(multi22[1][i22]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j22+0][i22+2]), .Out(multi22[2][i22]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j22+0][i22+3]), .Out(multi22[3][i22]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j22+0][i22+4]), .Out(multi22[4][i22]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j22+1][i22+0]), .Out(multi22[5][i22]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j22+1][i22+1]), .Out(multi22[6][i22]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j22+1][i22+2]), .Out(multi22[7][i22]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j22+1][i22+3]), .Out(multi22[8][i22]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j22+1][i22+4]), .Out(multi22[9][i22]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j22+2][i22+0]), .Out(multi22[10][i22]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j22+2][i22+1]), .Out(multi22[11][i22]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j22+2][i22+2]), .Out(multi22[12][i22]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j22+2][i22+3]), .Out(multi22[13][i22]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j22+2][i22+4]), .Out(multi22[14][i22]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j22+3][i22+0]), .Out(multi22[15][i22]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j22+3][i22+1]), .Out(multi22[16][i22]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j22+3][i22+2]), .Out(multi22[17][i22]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j22+3][i22+3]), .Out(multi22[18][i22]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j22+3][i22+4]), .Out(multi22[19][i22]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j22+4][i22+0]), .Out(multi22[20][i22]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j22+4][i22+1]), .Out(multi22[21][i22]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j22+4][i22+2]), .Out(multi22[22][i22]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j22+4][i22+3]), .Out(multi22[23][i22]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j22+4][i22+4]), .Out(multi22[24][i22]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi22[0][i22]), .B(multi22[1][i22]), .Out(sum22[0][i22]));
      FP16_Add stage026(.A(multi22[2][i22]), .B(multi22[3][i22]), .Out(sum22[1][i22]));
      FP16_Add stage027(.A(multi22[4][i22]), .B(multi22[5][i22]), .Out(sum22[2][i22]));
      FP16_Add stage028(.A(multi22[6][i22]), .B(multi22[7][i22]), .Out(sum22[3][i22]));
      FP16_Add stage029(.A(multi22[8][i22]), .B(multi22[9][i22]), .Out(sum22[4][i22]));
      FP16_Add stage030(.A(multi22[10][i22]), .B(multi22[11][i22]), .Out(sum22[5][i22]));
      FP16_Add stage031(.A(multi22[12][i22]), .B(multi22[13][i22]), .Out(sum22[6][i22]));
      FP16_Add stage032(.A(multi22[14][i22]), .B(multi22[15][i22]), .Out(sum22[7][i22]));
      FP16_Add stage033(.A(multi22[16][i22]), .B(multi22[17][i22]), .Out(sum22[8][i22]));
      FP16_Add stage034(.A(multi22[18][i22]), .B(multi22[19][i22]), .Out(sum22[9][i22]));
      FP16_Add stage035(.A(multi22[20][i22]), .B(multi22[21][i22]), .Out(sum22[10][i22]));
      FP16_Add stage036(.A(multi22[22][i22]), .B(multi22[23][i22]), .Out(sum22[11][i22]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum22[0][i22]), .B(sum22[1][i22]), .Out(sum22[12][i22]));
      FP16_Add stage038(.A(sum22[2][i22]), .B(sum22[3][i22]), .Out(sum22[13][i22]));
      FP16_Add stage039(.A(sum22[4][i22]), .B(sum22[5][i22]), .Out(sum22[14][i22]));
      FP16_Add stage040(.A(sum22[6][i22]), .B(sum22[7][i22]), .Out(sum22[15][i22]));
      FP16_Add stage041(.A(sum22[8][i22]), .B(sum22[9][i22]), .Out(sum22[16][i22]));
      FP16_Add stage042(.A(sum22[10][i22]), .B(sum22[11][i22]), .Out(sum22[17][i22]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum22[12][i22]), .B(sum22[13][i22]), .Out(sum22[18][i22]));
      FP16_Add stage044(.A(sum22[14][i22]), .B(sum22[15][i22]), .Out(sum22[19][i22]));
      FP16_Add stage045(.A(sum22[16][i22]), .B(sum22[17][i22]), .Out(sum22[20][i22]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum22[18][i22]), .B(sum22[19][i22]), .Out(sum22[21][i22]));
      FP16_Add stage047(.A(sum22[20][i22]), .B(multi22[24][i22]), .Out(sum22[22][i22]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum22[21][i22]), .B(sum22[22][i22]), .Out(sum22[23][i22]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum22[23][i22]), .B(feature1Bias), .Out(data_11_array[j22][i22]));
    end
  endgenerate

////ROW 23
  generate
    localparam integer j23 = 23;
    for (i23 = 0; i23 < 24; i23 = i23 + 1)
    begin: addbit23
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature1Weight_0), .B(data_array[j23+0][i23+0]), .Out(multi23[0][i23]));
      FP16_Multiply stage01(.A(feature1Weight_1), .B(data_array[j23+0][i23+1]), .Out(multi23[1][i23]));
      FP16_Multiply stage02(.A(feature1Weight_2), .B(data_array[j23+0][i23+2]), .Out(multi23[2][i23]));
      FP16_Multiply stage03(.A(feature1Weight_3), .B(data_array[j23+0][i23+3]), .Out(multi23[3][i23]));
      FP16_Multiply stage04(.A(feature1Weight_4), .B(data_array[j23+0][i23+4]), .Out(multi23[4][i23]));
      FP16_Multiply stage05(.A(feature1Weight_5), .B(data_array[j23+1][i23+0]), .Out(multi23[5][i23]));
      FP16_Multiply stage06(.A(feature1Weight_6), .B(data_array[j23+1][i23+1]), .Out(multi23[6][i23]));
      FP16_Multiply stage07(.A(feature1Weight_7), .B(data_array[j23+1][i23+2]), .Out(multi23[7][i23]));
      FP16_Multiply stage08(.A(feature1Weight_8), .B(data_array[j23+1][i23+3]), .Out(multi23[8][i23]));
      FP16_Multiply stage09(.A(feature1Weight_9), .B(data_array[j23+1][i23+4]), .Out(multi23[9][i23]));
      FP16_Multiply stage010(.A(feature1Weight_10), .B(data_array[j23+2][i23+0]), .Out(multi23[10][i23]));
      FP16_Multiply stage011(.A(feature1Weight_11), .B(data_array[j23+2][i23+1]), .Out(multi23[11][i23]));
      FP16_Multiply stage012(.A(feature1Weight_12), .B(data_array[j23+2][i23+2]), .Out(multi23[12][i23]));
      FP16_Multiply stage013(.A(feature1Weight_13), .B(data_array[j23+2][i23+3]), .Out(multi23[13][i23]));
      FP16_Multiply stage014(.A(feature1Weight_14), .B(data_array[j23+2][i23+4]), .Out(multi23[14][i23]));
      FP16_Multiply stage015(.A(feature1Weight_15), .B(data_array[j23+3][i23+0]), .Out(multi23[15][i23]));
      FP16_Multiply stage016(.A(feature1Weight_16), .B(data_array[j23+3][i23+1]), .Out(multi23[16][i23]));
      FP16_Multiply stage017(.A(feature1Weight_17), .B(data_array[j23+3][i23+2]), .Out(multi23[17][i23]));
      FP16_Multiply stage018(.A(feature1Weight_18), .B(data_array[j23+3][i23+3]), .Out(multi23[18][i23]));
      FP16_Multiply stage019(.A(feature1Weight_19), .B(data_array[j23+3][i23+4]), .Out(multi23[19][i23]));
      FP16_Multiply stage020(.A(feature1Weight_20), .B(data_array[j23+4][i23+0]), .Out(multi23[20][i23]));
      FP16_Multiply stage021(.A(feature1Weight_21), .B(data_array[j23+4][i23+1]), .Out(multi23[21][i23]));
      FP16_Multiply stage022(.A(feature1Weight_22), .B(data_array[j23+4][i23+2]), .Out(multi23[22][i23]));
      FP16_Multiply stage023(.A(feature1Weight_23), .B(data_array[j23+4][i23+3]), .Out(multi23[23][i23]));
      FP16_Multiply stage024(.A(feature1Weight_24), .B(data_array[j23+4][i23+4]), .Out(multi23[24][i23]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi23[0][i23]), .B(multi23[1][i23]), .Out(sum23[0][i23]));
      FP16_Add stage026(.A(multi23[2][i23]), .B(multi23[3][i23]), .Out(sum23[1][i23]));
      FP16_Add stage027(.A(multi23[4][i23]), .B(multi23[5][i23]), .Out(sum23[2][i23]));
      FP16_Add stage028(.A(multi23[6][i23]), .B(multi23[7][i23]), .Out(sum23[3][i23]));
      FP16_Add stage029(.A(multi23[8][i23]), .B(multi23[9][i23]), .Out(sum23[4][i23]));
      FP16_Add stage030(.A(multi23[10][i23]), .B(multi23[11][i23]), .Out(sum23[5][i23]));
      FP16_Add stage031(.A(multi23[12][i23]), .B(multi23[13][i23]), .Out(sum23[6][i23]));
      FP16_Add stage032(.A(multi23[14][i23]), .B(multi23[15][i23]), .Out(sum23[7][i23]));
      FP16_Add stage033(.A(multi23[16][i23]), .B(multi23[17][i23]), .Out(sum23[8][i23]));
      FP16_Add stage034(.A(multi23[18][i23]), .B(multi23[19][i23]), .Out(sum23[9][i23]));
      FP16_Add stage035(.A(multi23[20][i23]), .B(multi23[21][i23]), .Out(sum23[10][i23]));
      FP16_Add stage036(.A(multi23[22][i23]), .B(multi23[23][i23]), .Out(sum23[11][i23]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum23[0][i23]), .B(sum23[1][i23]), .Out(sum23[12][i23]));
      FP16_Add stage038(.A(sum23[2][i23]), .B(sum23[3][i23]), .Out(sum23[13][i23]));
      FP16_Add stage039(.A(sum23[4][i23]), .B(sum23[5][i23]), .Out(sum23[14][i23]));
      FP16_Add stage040(.A(sum23[6][i23]), .B(sum23[7][i23]), .Out(sum23[15][i23]));
      FP16_Add stage041(.A(sum23[8][i23]), .B(sum23[9][i23]), .Out(sum23[16][i23]));
      FP16_Add stage042(.A(sum23[10][i23]), .B(sum23[11][i23]), .Out(sum23[17][i23]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum23[12][i23]), .B(sum23[13][i23]), .Out(sum23[18][i23]));
      FP16_Add stage044(.A(sum23[14][i23]), .B(sum23[15][i23]), .Out(sum23[19][i23]));
      FP16_Add stage045(.A(sum23[16][i23]), .B(sum23[17][i23]), .Out(sum23[20][i23]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum23[18][i23]), .B(sum23[19][i23]), .Out(sum23[21][i23]));
      FP16_Add stage047(.A(sum23[20][i23]), .B(multi23[24][i23]), .Out(sum23[22][i23]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum23[21][i23]), .B(sum23[22][i23]), .Out(sum23[23][i23]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum23[23][i23]), .B(feature1Bias), .Out(data_11_array[j23][i23]));
    end
  endgenerate
  
  localparam integer c0 = 0;
    generate 
        localparam integer d0 = 0;
        for (n0 = 0; n0 < 16; n0 = n0 + 1) 
        begin: outbit0
            assign data_11[n0 + d0*16 + c0*28*16] = data_11_array[c0][d0][n0];
        end
    endgenerate
    generate 
        localparam integer d1 = 1;
        for (n1 = 0; n1 < 16; n1 = n1 + 1) 
        begin: outbit1
            assign data_11[n1 + d1*16 + c0*28*16] = data_11_array[c0][d1][n1];
        end
    endgenerate
    generate 
        localparam integer d2 = 2;
        for (n2 = 0; n2 < 16; n2 = n2 + 1) 
        begin: outbit2
            assign data_11[n2 + d2*16 + c0*28*16] = data_11_array[c0][d2][n2];
        end
    endgenerate
    generate 
        localparam integer d3 = 3;
        for (n3 = 0; n3 < 16; n3 = n3 + 1) 
        begin: outbit3
            assign data_11[n3 + d3*16 + c0*28*16] = data_11_array[c0][d3][n3];
        end
    endgenerate
    generate 
        localparam integer d4 = 4;
        for (n4 = 0; n4 < 16; n4 = n4 + 1) 
        begin: outbit4
            assign data_11[n4 + d4*16 + c0*28*16] = data_11_array[c0][d4][n4];
        end
    endgenerate
    generate 
        localparam integer d5 = 5;
        for (n5 = 0; n5 < 16; n5 = n5 + 1) 
        begin: outbit5
            assign data_11[n5 + d5*16 + c0*28*16] = data_11_array[c0][d5][n5];
        end
    endgenerate
    generate 
        localparam integer d6 = 6;
        for (n6 = 0; n6 < 16; n6 = n6 + 1) 
        begin: outbit6
            assign data_11[n6 + d6*16 + c0*28*16] = data_11_array[c0][d6][n6];
        end
    endgenerate
    generate 
        localparam integer d7 = 7;
        for (n7 = 0; n7 < 16; n7 = n7 + 1) 
        begin: outbit7
            assign data_11[n7 + d7*16 + c0*28*16] = data_11_array[c0][d7][n7];
        end
    endgenerate
    generate 
        localparam integer d8 = 8;
        for (n8 = 0; n8 < 16; n8 = n8 + 1) 
        begin: outbit8
            assign data_11[n8 + d8*16 + c0*28*16] = data_11_array[c0][d8][n8];
        end
    endgenerate
    generate 
        localparam integer d9 = 9;
        for (n9 = 0; n9 < 16; n9 = n9 + 1) 
        begin: outbit9
            assign data_11[n9 + d9*16 + c0*28*16] = data_11_array[c0][d9][n9];
        end
    endgenerate
    generate 
        localparam integer d10 = 10;
        for (n10 = 0; n10 < 16; n10 = n10 + 1) 
        begin: outbit10
            assign data_11[n10 + d10*16 + c0*28*16] = data_11_array[c0][d10][n10];
        end
    endgenerate
    generate 
        localparam integer d11 = 11;
        for (n11 = 0; n11 < 16; n11 = n11 + 1) 
        begin: outbit11
            assign data_11[n11 + d11*16 + c0*28*16] = data_11_array[c0][d11][n11];
        end
    endgenerate
    generate 
        localparam integer d12 = 12;
        for (n12 = 0; n12 < 16; n12 = n12 + 1) 
        begin: outbit12
            assign data_11[n12 + d12*16 + c0*28*16] = data_11_array[c0][d12][n12];
        end
    endgenerate
    generate 
        localparam integer d13 = 13;
        for (n13 = 0; n13 < 16; n13 = n13 + 1) 
        begin: outbit13
            assign data_11[n13 + d13*16 + c0*28*16] = data_11_array[c0][d13][n13];
        end
    endgenerate
    generate 
        localparam integer d14 = 14;
        for (n14 = 0; n14 < 16; n14 = n14 + 1) 
        begin: outbit14
            assign data_11[n14 + d14*16 + c0*28*16] = data_11_array[c0][d14][n14];
        end
    endgenerate
    generate 
        localparam integer d15 = 15;
        for (n15 = 0; n15 < 16; n15 = n15 + 1) 
        begin: outbit15
            assign data_11[n15 + d15*16 + c0*28*16] = data_11_array[c0][d15][n15];
        end
    endgenerate
    generate 
        localparam integer d16 = 16;
        for (n16 = 0; n16 < 16; n16 = n16 + 1) 
        begin: outbit16
            assign data_11[n16 + d16*16 + c0*28*16] = data_11_array[c0][d16][n16];
        end
    endgenerate
    generate 
        localparam integer d17 = 17;
        for (n17 = 0; n17 < 16; n17 = n17 + 1) 
        begin: outbit17
            assign data_11[n17 + d17*16 + c0*28*16] = data_11_array[c0][d17][n17];
        end
    endgenerate
    generate 
        localparam integer d18 = 18;
        for (n18 = 0; n18 < 16; n18 = n18 + 1) 
        begin: outbit18
            assign data_11[n18 + d18*16 + c0*28*16] = data_11_array[c0][d18][n18];
        end
    endgenerate
    generate 
        localparam integer d19 = 19;
        for (n19 = 0; n19 < 16; n19 = n19 + 1) 
        begin: outbit19
            assign data_11[n19 + d19*16 + c0*28*16] = data_11_array[c0][d19][n19];
        end
    endgenerate
    generate 
        localparam integer d20 = 20;
        for (n20 = 0; n20 < 16; n20 = n20 + 1) 
        begin: outbit20
            assign data_11[n20 + d20*16 + c0*28*16] = data_11_array[c0][d20][n20];
        end
    endgenerate
    generate 
        localparam integer d21 = 21;
        for (n21 = 0; n21 < 16; n21 = n21 + 1) 
        begin: outbit21
            assign data_11[n21 + d21*16 + c0*28*16] = data_11_array[c0][d21][n21];
        end
    endgenerate
    generate 
        localparam integer d22 = 22;
        for (n22 = 0; n22 < 16; n22 = n22 + 1) 
        begin: outbit22
            assign data_11[n22 + d22*16 + c0*28*16] = data_11_array[c0][d22][n22];
        end
    endgenerate
    generate 
        localparam integer d23 = 23;
        for (n23 = 0; n23 < 16; n23 = n23 + 1) 
        begin: outbit23
            assign data_11[n23 + d23*16 + c0*28*16] = data_11_array[c0][d23][n23];
        end
    endgenerate
    generate 
        localparam integer d24 = 24;
        for (n24 = 0; n24 < 16; n24 = n24 + 1) 
        begin: outbit24
            assign data_11[n24 + d24*16 + c0*28*16] = data_11_array[c0][d24][n24];
        end
    endgenerate
    generate 
        localparam integer d25 = 25;
        for (n25 = 0; n25 < 16; n25 = n25 + 1) 
        begin: outbit25
            assign data_11[n25 + d25*16 + c0*28*16] = data_11_array[c0][d25][n25];
        end
    endgenerate
    generate 
        localparam integer d26 = 26;
        for (n26 = 0; n26 < 16; n26 = n26 + 1) 
        begin: outbit26
            assign data_11[n26 + d26*16 + c0*28*16] = data_11_array[c0][d26][n26];
        end
    endgenerate
    generate 
        localparam integer d27 = 27;
        for (n27 = 0; n27 < 16; n27 = n27 + 1) 
        begin: outbit27
            assign data_11[n27 + d27*16 + c0*28*16] = data_11_array[c0][d27][n27];
        end
    endgenerate
    localparam integer c1 = 1;
    generate 
        localparam integer d28 = 0;
        for (n28 = 0; n28 < 16; n28 = n28 + 1) 
        begin: outbit28
            assign data_11[n28 + d28*16 + c1*28*16] = data_11_array[c1][d28][n28];
        end
    endgenerate
    generate 
        localparam integer d29 = 1;
        for (n29 = 0; n29 < 16; n29 = n29 + 1) 
        begin: outbit29
            assign data_11[n29 + d29*16 + c1*28*16] = data_11_array[c1][d29][n29];
        end
    endgenerate
    generate 
        localparam integer d30 = 2;
        for (n30 = 0; n30 < 16; n30 = n30 + 1) 
        begin: outbit30
            assign data_11[n30 + d30*16 + c1*28*16] = data_11_array[c1][d30][n30];
        end
    endgenerate
    generate 
        localparam integer d31 = 3;
        for (n31 = 0; n31 < 16; n31 = n31 + 1) 
        begin: outbit31
            assign data_11[n31 + d31*16 + c1*28*16] = data_11_array[c1][d31][n31];
        end
    endgenerate
    generate 
        localparam integer d32 = 4;
        for (n32 = 0; n32 < 16; n32 = n32 + 1) 
        begin: outbit32
            assign data_11[n32 + d32*16 + c1*28*16] = data_11_array[c1][d32][n32];
        end
    endgenerate
    generate 
        localparam integer d33 = 5;
        for (n33 = 0; n33 < 16; n33 = n33 + 1) 
        begin: outbit33
            assign data_11[n33 + d33*16 + c1*28*16] = data_11_array[c1][d33][n33];
        end
    endgenerate
    generate 
        localparam integer d34 = 6;
        for (n34 = 0; n34 < 16; n34 = n34 + 1) 
        begin: outbit34
            assign data_11[n34 + d34*16 + c1*28*16] = data_11_array[c1][d34][n34];
        end
    endgenerate
    generate 
        localparam integer d35 = 7;
        for (n35 = 0; n35 < 16; n35 = n35 + 1) 
        begin: outbit35
            assign data_11[n35 + d35*16 + c1*28*16] = data_11_array[c1][d35][n35];
        end
    endgenerate
    generate 
        localparam integer d36 = 8;
        for (n36 = 0; n36 < 16; n36 = n36 + 1) 
        begin: outbit36
            assign data_11[n36 + d36*16 + c1*28*16] = data_11_array[c1][d36][n36];
        end
    endgenerate
    generate 
        localparam integer d37 = 9;
        for (n37 = 0; n37 < 16; n37 = n37 + 1) 
        begin: outbit37
            assign data_11[n37 + d37*16 + c1*28*16] = data_11_array[c1][d37][n37];
        end
    endgenerate
    generate 
        localparam integer d38 = 10;
        for (n38 = 0; n38 < 16; n38 = n38 + 1) 
        begin: outbit38
            assign data_11[n38 + d38*16 + c1*28*16] = data_11_array[c1][d38][n38];
        end
    endgenerate
    generate 
        localparam integer d39 = 11;
        for (n39 = 0; n39 < 16; n39 = n39 + 1) 
        begin: outbit39
            assign data_11[n39 + d39*16 + c1*28*16] = data_11_array[c1][d39][n39];
        end
    endgenerate
    generate 
        localparam integer d40 = 12;
        for (n40 = 0; n40 < 16; n40 = n40 + 1) 
        begin: outbit40
            assign data_11[n40 + d40*16 + c1*28*16] = data_11_array[c1][d40][n40];
        end
    endgenerate
    generate 
        localparam integer d41 = 13;
        for (n41 = 0; n41 < 16; n41 = n41 + 1) 
        begin: outbit41
            assign data_11[n41 + d41*16 + c1*28*16] = data_11_array[c1][d41][n41];
        end
    endgenerate
    generate 
        localparam integer d42 = 14;
        for (n42 = 0; n42 < 16; n42 = n42 + 1) 
        begin: outbit42
            assign data_11[n42 + d42*16 + c1*28*16] = data_11_array[c1][d42][n42];
        end
    endgenerate
    generate 
        localparam integer d43 = 15;
        for (n43 = 0; n43 < 16; n43 = n43 + 1) 
        begin: outbit43
            assign data_11[n43 + d43*16 + c1*28*16] = data_11_array[c1][d43][n43];
        end
    endgenerate
    generate 
        localparam integer d44 = 16;
        for (n44 = 0; n44 < 16; n44 = n44 + 1) 
        begin: outbit44
            assign data_11[n44 + d44*16 + c1*28*16] = data_11_array[c1][d44][n44];
        end
    endgenerate
    generate 
        localparam integer d45 = 17;
        for (n45 = 0; n45 < 16; n45 = n45 + 1) 
        begin: outbit45
            assign data_11[n45 + d45*16 + c1*28*16] = data_11_array[c1][d45][n45];
        end
    endgenerate
    generate 
        localparam integer d46 = 18;
        for (n46 = 0; n46 < 16; n46 = n46 + 1) 
        begin: outbit46
            assign data_11[n46 + d46*16 + c1*28*16] = data_11_array[c1][d46][n46];
        end
    endgenerate
    generate 
        localparam integer d47 = 19;
        for (n47 = 0; n47 < 16; n47 = n47 + 1) 
        begin: outbit47
            assign data_11[n47 + d47*16 + c1*28*16] = data_11_array[c1][d47][n47];
        end
    endgenerate
    generate 
        localparam integer d48 = 20;
        for (n48 = 0; n48 < 16; n48 = n48 + 1) 
        begin: outbit48
            assign data_11[n48 + d48*16 + c1*28*16] = data_11_array[c1][d48][n48];
        end
    endgenerate
    generate 
        localparam integer d49 = 21;
        for (n49 = 0; n49 < 16; n49 = n49 + 1) 
        begin: outbit49
            assign data_11[n49 + d49*16 + c1*28*16] = data_11_array[c1][d49][n49];
        end
    endgenerate
    generate 
        localparam integer d50 = 22;
        for (n50 = 0; n50 < 16; n50 = n50 + 1) 
        begin: outbit50
            assign data_11[n50 + d50*16 + c1*28*16] = data_11_array[c1][d50][n50];
        end
    endgenerate
    generate 
        localparam integer d51 = 23;
        for (n51 = 0; n51 < 16; n51 = n51 + 1) 
        begin: outbit51
            assign data_11[n51 + d51*16 + c1*28*16] = data_11_array[c1][d51][n51];
        end
    endgenerate
    generate 
        localparam integer d52 = 24;
        for (n52 = 0; n52 < 16; n52 = n52 + 1) 
        begin: outbit52
            assign data_11[n52 + d52*16 + c1*28*16] = data_11_array[c1][d52][n52];
        end
    endgenerate
    generate 
        localparam integer d53 = 25;
        for (n53 = 0; n53 < 16; n53 = n53 + 1) 
        begin: outbit53
            assign data_11[n53 + d53*16 + c1*28*16] = data_11_array[c1][d53][n53];
        end
    endgenerate
    generate 
        localparam integer d54 = 26;
        for (n54 = 0; n54 < 16; n54 = n54 + 1) 
        begin: outbit54
            assign data_11[n54 + d54*16 + c1*28*16] = data_11_array[c1][d54][n54];
        end
    endgenerate
    generate 
        localparam integer d55 = 27;
        for (n55 = 0; n55 < 16; n55 = n55 + 1) 
        begin: outbit55
            assign data_11[n55 + d55*16 + c1*28*16] = data_11_array[c1][d55][n55];
        end
    endgenerate
    localparam integer c2 = 2;
    generate 
        localparam integer d56 = 0;
        for (n56 = 0; n56 < 16; n56 = n56 + 1) 
        begin: outbit56
            assign data_11[n56 + d56*16 + c2*28*16] = data_11_array[c2][d56][n56];
        end
    endgenerate
    generate 
        localparam integer d57 = 1;
        for (n57 = 0; n57 < 16; n57 = n57 + 1) 
        begin: outbit57
            assign data_11[n57 + d57*16 + c2*28*16] = data_11_array[c2][d57][n57];
        end
    endgenerate
    generate 
        localparam integer d58 = 2;
        for (n58 = 0; n58 < 16; n58 = n58 + 1) 
        begin: outbit58
            assign data_11[n58 + d58*16 + c2*28*16] = data_11_array[c2][d58][n58];
        end
    endgenerate
    generate 
        localparam integer d59 = 3;
        for (n59 = 0; n59 < 16; n59 = n59 + 1) 
        begin: outbit59
            assign data_11[n59 + d59*16 + c2*28*16] = data_11_array[c2][d59][n59];
        end
    endgenerate
    generate 
        localparam integer d60 = 4;
        for (n60 = 0; n60 < 16; n60 = n60 + 1) 
        begin: outbit60
            assign data_11[n60 + d60*16 + c2*28*16] = data_11_array[c2][d60][n60];
        end
    endgenerate
    generate 
        localparam integer d61 = 5;
        for (n61 = 0; n61 < 16; n61 = n61 + 1) 
        begin: outbit61
            assign data_11[n61 + d61*16 + c2*28*16] = data_11_array[c2][d61][n61];
        end
    endgenerate
    generate 
        localparam integer d62 = 6;
        for (n62 = 0; n62 < 16; n62 = n62 + 1) 
        begin: outbit62
            assign data_11[n62 + d62*16 + c2*28*16] = data_11_array[c2][d62][n62];
        end
    endgenerate
    generate 
        localparam integer d63 = 7;
        for (n63 = 0; n63 < 16; n63 = n63 + 1) 
        begin: outbit63
            assign data_11[n63 + d63*16 + c2*28*16] = data_11_array[c2][d63][n63];
        end
    endgenerate
    generate 
        localparam integer d64 = 8;
        for (n64 = 0; n64 < 16; n64 = n64 + 1) 
        begin: outbit64
            assign data_11[n64 + d64*16 + c2*28*16] = data_11_array[c2][d64][n64];
        end
    endgenerate
    generate 
        localparam integer d65 = 9;
        for (n65 = 0; n65 < 16; n65 = n65 + 1) 
        begin: outbit65
            assign data_11[n65 + d65*16 + c2*28*16] = data_11_array[c2][d65][n65];
        end
    endgenerate
    generate 
        localparam integer d66 = 10;
        for (n66 = 0; n66 < 16; n66 = n66 + 1) 
        begin: outbit66
            assign data_11[n66 + d66*16 + c2*28*16] = data_11_array[c2][d66][n66];
        end
    endgenerate
    generate 
        localparam integer d67 = 11;
        for (n67 = 0; n67 < 16; n67 = n67 + 1) 
        begin: outbit67
            assign data_11[n67 + d67*16 + c2*28*16] = data_11_array[c2][d67][n67];
        end
    endgenerate
    generate 
        localparam integer d68 = 12;
        for (n68 = 0; n68 < 16; n68 = n68 + 1) 
        begin: outbit68
            assign data_11[n68 + d68*16 + c2*28*16] = data_11_array[c2][d68][n68];
        end
    endgenerate
    generate 
        localparam integer d69 = 13;
        for (n69 = 0; n69 < 16; n69 = n69 + 1) 
        begin: outbit69
            assign data_11[n69 + d69*16 + c2*28*16] = data_11_array[c2][d69][n69];
        end
    endgenerate
    generate 
        localparam integer d70 = 14;
        for (n70 = 0; n70 < 16; n70 = n70 + 1) 
        begin: outbit70
            assign data_11[n70 + d70*16 + c2*28*16] = data_11_array[c2][d70][n70];
        end
    endgenerate
    generate 
        localparam integer d71 = 15;
        for (n71 = 0; n71 < 16; n71 = n71 + 1) 
        begin: outbit71
            assign data_11[n71 + d71*16 + c2*28*16] = data_11_array[c2][d71][n71];
        end
    endgenerate
    generate 
        localparam integer d72 = 16;
        for (n72 = 0; n72 < 16; n72 = n72 + 1) 
        begin: outbit72
            assign data_11[n72 + d72*16 + c2*28*16] = data_11_array[c2][d72][n72];
        end
    endgenerate
    generate 
        localparam integer d73 = 17;
        for (n73 = 0; n73 < 16; n73 = n73 + 1) 
        begin: outbit73
            assign data_11[n73 + d73*16 + c2*28*16] = data_11_array[c2][d73][n73];
        end
    endgenerate
    generate 
        localparam integer d74 = 18;
        for (n74 = 0; n74 < 16; n74 = n74 + 1) 
        begin: outbit74
            assign data_11[n74 + d74*16 + c2*28*16] = data_11_array[c2][d74][n74];
        end
    endgenerate
    generate 
        localparam integer d75 = 19;
        for (n75 = 0; n75 < 16; n75 = n75 + 1) 
        begin: outbit75
            assign data_11[n75 + d75*16 + c2*28*16] = data_11_array[c2][d75][n75];
        end
    endgenerate
    generate 
        localparam integer d76 = 20;
        for (n76 = 0; n76 < 16; n76 = n76 + 1) 
        begin: outbit76
            assign data_11[n76 + d76*16 + c2*28*16] = data_11_array[c2][d76][n76];
        end
    endgenerate
    generate 
        localparam integer d77 = 21;
        for (n77 = 0; n77 < 16; n77 = n77 + 1) 
        begin: outbit77
            assign data_11[n77 + d77*16 + c2*28*16] = data_11_array[c2][d77][n77];
        end
    endgenerate
    generate 
        localparam integer d78 = 22;
        for (n78 = 0; n78 < 16; n78 = n78 + 1) 
        begin: outbit78
            assign data_11[n78 + d78*16 + c2*28*16] = data_11_array[c2][d78][n78];
        end
    endgenerate
    generate 
        localparam integer d79 = 23;
        for (n79 = 0; n79 < 16; n79 = n79 + 1) 
        begin: outbit79
            assign data_11[n79 + d79*16 + c2*28*16] = data_11_array[c2][d79][n79];
        end
    endgenerate
    generate 
        localparam integer d80 = 24;
        for (n80 = 0; n80 < 16; n80 = n80 + 1) 
        begin: outbit80
            assign data_11[n80 + d80*16 + c2*28*16] = data_11_array[c2][d80][n80];
        end
    endgenerate
    generate 
        localparam integer d81 = 25;
        for (n81 = 0; n81 < 16; n81 = n81 + 1) 
        begin: outbit81
            assign data_11[n81 + d81*16 + c2*28*16] = data_11_array[c2][d81][n81];
        end
    endgenerate
    generate 
        localparam integer d82 = 26;
        for (n82 = 0; n82 < 16; n82 = n82 + 1) 
        begin: outbit82
            assign data_11[n82 + d82*16 + c2*28*16] = data_11_array[c2][d82][n82];
        end
    endgenerate
    generate 
        localparam integer d83 = 27;
        for (n83 = 0; n83 < 16; n83 = n83 + 1) 
        begin: outbit83
            assign data_11[n83 + d83*16 + c2*28*16] = data_11_array[c2][d83][n83];
        end
    endgenerate
    localparam integer c3 = 3;
    generate 
        localparam integer d84 = 0;
        for (n84 = 0; n84 < 16; n84 = n84 + 1) 
        begin: outbit84
            assign data_11[n84 + d84*16 + c3*28*16] = data_11_array[c3][d84][n84];
        end
    endgenerate
    generate 
        localparam integer d85 = 1;
        for (n85 = 0; n85 < 16; n85 = n85 + 1) 
        begin: outbit85
            assign data_11[n85 + d85*16 + c3*28*16] = data_11_array[c3][d85][n85];
        end
    endgenerate
    generate 
        localparam integer d86 = 2;
        for (n86 = 0; n86 < 16; n86 = n86 + 1) 
        begin: outbit86
            assign data_11[n86 + d86*16 + c3*28*16] = data_11_array[c3][d86][n86];
        end
    endgenerate
    generate 
        localparam integer d87 = 3;
        for (n87 = 0; n87 < 16; n87 = n87 + 1) 
        begin: outbit87
            assign data_11[n87 + d87*16 + c3*28*16] = data_11_array[c3][d87][n87];
        end
    endgenerate
    generate 
        localparam integer d88 = 4;
        for (n88 = 0; n88 < 16; n88 = n88 + 1) 
        begin: outbit88
            assign data_11[n88 + d88*16 + c3*28*16] = data_11_array[c3][d88][n88];
        end
    endgenerate
    generate 
        localparam integer d89 = 5;
        for (n89 = 0; n89 < 16; n89 = n89 + 1) 
        begin: outbit89
            assign data_11[n89 + d89*16 + c3*28*16] = data_11_array[c3][d89][n89];
        end
    endgenerate
    generate 
        localparam integer d90 = 6;
        for (n90 = 0; n90 < 16; n90 = n90 + 1) 
        begin: outbit90
            assign data_11[n90 + d90*16 + c3*28*16] = data_11_array[c3][d90][n90];
        end
    endgenerate
    generate 
        localparam integer d91 = 7;
        for (n91 = 0; n91 < 16; n91 = n91 + 1) 
        begin: outbit91
            assign data_11[n91 + d91*16 + c3*28*16] = data_11_array[c3][d91][n91];
        end
    endgenerate
    generate 
        localparam integer d92 = 8;
        for (n92 = 0; n92 < 16; n92 = n92 + 1) 
        begin: outbit92
            assign data_11[n92 + d92*16 + c3*28*16] = data_11_array[c3][d92][n92];
        end
    endgenerate
    generate 
        localparam integer d93 = 9;
        for (n93 = 0; n93 < 16; n93 = n93 + 1) 
        begin: outbit93
            assign data_11[n93 + d93*16 + c3*28*16] = data_11_array[c3][d93][n93];
        end
    endgenerate
    generate 
        localparam integer d94 = 10;
        for (n94 = 0; n94 < 16; n94 = n94 + 1) 
        begin: outbit94
            assign data_11[n94 + d94*16 + c3*28*16] = data_11_array[c3][d94][n94];
        end
    endgenerate
    generate 
        localparam integer d95 = 11;
        for (n95 = 0; n95 < 16; n95 = n95 + 1) 
        begin: outbit95
            assign data_11[n95 + d95*16 + c3*28*16] = data_11_array[c3][d95][n95];
        end
    endgenerate
    generate 
        localparam integer d96 = 12;
        for (n96 = 0; n96 < 16; n96 = n96 + 1) 
        begin: outbit96
            assign data_11[n96 + d96*16 + c3*28*16] = data_11_array[c3][d96][n96];
        end
    endgenerate
    generate 
        localparam integer d97 = 13;
        for (n97 = 0; n97 < 16; n97 = n97 + 1) 
        begin: outbit97
            assign data_11[n97 + d97*16 + c3*28*16] = data_11_array[c3][d97][n97];
        end
    endgenerate
    generate 
        localparam integer d98 = 14;
        for (n98 = 0; n98 < 16; n98 = n98 + 1) 
        begin: outbit98
            assign data_11[n98 + d98*16 + c3*28*16] = data_11_array[c3][d98][n98];
        end
    endgenerate
    generate 
        localparam integer d99 = 15;
        for (n99 = 0; n99 < 16; n99 = n99 + 1) 
        begin: outbit99
            assign data_11[n99 + d99*16 + c3*28*16] = data_11_array[c3][d99][n99];
        end
    endgenerate
    generate 
        localparam integer d100 = 16;
        for (n100 = 0; n100 < 16; n100 = n100 + 1) 
        begin: outbit100
            assign data_11[n100 + d100*16 + c3*28*16] = data_11_array[c3][d100][n100];
        end
    endgenerate
    generate 
        localparam integer d101 = 17;
        for (n101 = 0; n101 < 16; n101 = n101 + 1) 
        begin: outbit101
            assign data_11[n101 + d101*16 + c3*28*16] = data_11_array[c3][d101][n101];
        end
    endgenerate
    generate 
        localparam integer d102 = 18;
        for (n102 = 0; n102 < 16; n102 = n102 + 1) 
        begin: outbit102
            assign data_11[n102 + d102*16 + c3*28*16] = data_11_array[c3][d102][n102];
        end
    endgenerate
    generate 
        localparam integer d103 = 19;
        for (n103 = 0; n103 < 16; n103 = n103 + 1) 
        begin: outbit103
            assign data_11[n103 + d103*16 + c3*28*16] = data_11_array[c3][d103][n103];
        end
    endgenerate
    generate 
        localparam integer d104 = 20;
        for (n104 = 0; n104 < 16; n104 = n104 + 1) 
        begin: outbit104
            assign data_11[n104 + d104*16 + c3*28*16] = data_11_array[c3][d104][n104];
        end
    endgenerate
    generate 
        localparam integer d105 = 21;
        for (n105 = 0; n105 < 16; n105 = n105 + 1) 
        begin: outbit105
            assign data_11[n105 + d105*16 + c3*28*16] = data_11_array[c3][d105][n105];
        end
    endgenerate
    generate 
        localparam integer d106 = 22;
        for (n106 = 0; n106 < 16; n106 = n106 + 1) 
        begin: outbit106
            assign data_11[n106 + d106*16 + c3*28*16] = data_11_array[c3][d106][n106];
        end
    endgenerate
    generate 
        localparam integer d107 = 23;
        for (n107 = 0; n107 < 16; n107 = n107 + 1) 
        begin: outbit107
            assign data_11[n107 + d107*16 + c3*28*16] = data_11_array[c3][d107][n107];
        end
    endgenerate
    generate 
        localparam integer d108 = 24;
        for (n108 = 0; n108 < 16; n108 = n108 + 1) 
        begin: outbit108
            assign data_11[n108 + d108*16 + c3*28*16] = data_11_array[c3][d108][n108];
        end
    endgenerate
    generate 
        localparam integer d109 = 25;
        for (n109 = 0; n109 < 16; n109 = n109 + 1) 
        begin: outbit109
            assign data_11[n109 + d109*16 + c3*28*16] = data_11_array[c3][d109][n109];
        end
    endgenerate
    generate 
        localparam integer d110 = 26;
        for (n110 = 0; n110 < 16; n110 = n110 + 1) 
        begin: outbit110
            assign data_11[n110 + d110*16 + c3*28*16] = data_11_array[c3][d110][n110];
        end
    endgenerate
    generate 
        localparam integer d111 = 27;
        for (n111 = 0; n111 < 16; n111 = n111 + 1) 
        begin: outbit111
            assign data_11[n111 + d111*16 + c3*28*16] = data_11_array[c3][d111][n111];
        end
    endgenerate
    localparam integer c4 = 4;
    generate 
        localparam integer d112 = 0;
        for (n112 = 0; n112 < 16; n112 = n112 + 1) 
        begin: outbit112
            assign data_11[n112 + d112*16 + c4*28*16] = data_11_array[c4][d112][n112];
        end
    endgenerate
    generate 
        localparam integer d113 = 1;
        for (n113 = 0; n113 < 16; n113 = n113 + 1) 
        begin: outbit113
            assign data_11[n113 + d113*16 + c4*28*16] = data_11_array[c4][d113][n113];
        end
    endgenerate
    generate 
        localparam integer d114 = 2;
        for (n114 = 0; n114 < 16; n114 = n114 + 1) 
        begin: outbit114
            assign data_11[n114 + d114*16 + c4*28*16] = data_11_array[c4][d114][n114];
        end
    endgenerate
    generate 
        localparam integer d115 = 3;
        for (n115 = 0; n115 < 16; n115 = n115 + 1) 
        begin: outbit115
            assign data_11[n115 + d115*16 + c4*28*16] = data_11_array[c4][d115][n115];
        end
    endgenerate
    generate 
        localparam integer d116 = 4;
        for (n116 = 0; n116 < 16; n116 = n116 + 1) 
        begin: outbit116
            assign data_11[n116 + d116*16 + c4*28*16] = data_11_array[c4][d116][n116];
        end
    endgenerate
    generate 
        localparam integer d117 = 5;
        for (n117 = 0; n117 < 16; n117 = n117 + 1) 
        begin: outbit117
            assign data_11[n117 + d117*16 + c4*28*16] = data_11_array[c4][d117][n117];
        end
    endgenerate
    generate 
        localparam integer d118 = 6;
        for (n118 = 0; n118 < 16; n118 = n118 + 1) 
        begin: outbit118
            assign data_11[n118 + d118*16 + c4*28*16] = data_11_array[c4][d118][n118];
        end
    endgenerate
    generate 
        localparam integer d119 = 7;
        for (n119 = 0; n119 < 16; n119 = n119 + 1) 
        begin: outbit119
            assign data_11[n119 + d119*16 + c4*28*16] = data_11_array[c4][d119][n119];
        end
    endgenerate
    generate 
        localparam integer d120 = 8;
        for (n120 = 0; n120 < 16; n120 = n120 + 1) 
        begin: outbit120
            assign data_11[n120 + d120*16 + c4*28*16] = data_11_array[c4][d120][n120];
        end
    endgenerate
    generate 
        localparam integer d121 = 9;
        for (n121 = 0; n121 < 16; n121 = n121 + 1) 
        begin: outbit121
            assign data_11[n121 + d121*16 + c4*28*16] = data_11_array[c4][d121][n121];
        end
    endgenerate
    generate 
        localparam integer d122 = 10;
        for (n122 = 0; n122 < 16; n122 = n122 + 1) 
        begin: outbit122
            assign data_11[n122 + d122*16 + c4*28*16] = data_11_array[c4][d122][n122];
        end
    endgenerate
    generate 
        localparam integer d123 = 11;
        for (n123 = 0; n123 < 16; n123 = n123 + 1) 
        begin: outbit123
            assign data_11[n123 + d123*16 + c4*28*16] = data_11_array[c4][d123][n123];
        end
    endgenerate
    generate 
        localparam integer d124 = 12;
        for (n124 = 0; n124 < 16; n124 = n124 + 1) 
        begin: outbit124
            assign data_11[n124 + d124*16 + c4*28*16] = data_11_array[c4][d124][n124];
        end
    endgenerate
    generate 
        localparam integer d125 = 13;
        for (n125 = 0; n125 < 16; n125 = n125 + 1) 
        begin: outbit125
            assign data_11[n125 + d125*16 + c4*28*16] = data_11_array[c4][d125][n125];
        end
    endgenerate
    generate 
        localparam integer d126 = 14;
        for (n126 = 0; n126 < 16; n126 = n126 + 1) 
        begin: outbit126
            assign data_11[n126 + d126*16 + c4*28*16] = data_11_array[c4][d126][n126];
        end
    endgenerate
    generate 
        localparam integer d127 = 15;
        for (n127 = 0; n127 < 16; n127 = n127 + 1) 
        begin: outbit127
            assign data_11[n127 + d127*16 + c4*28*16] = data_11_array[c4][d127][n127];
        end
    endgenerate
    generate 
        localparam integer d128 = 16;
        for (n128 = 0; n128 < 16; n128 = n128 + 1) 
        begin: outbit128
            assign data_11[n128 + d128*16 + c4*28*16] = data_11_array[c4][d128][n128];
        end
    endgenerate
    generate 
        localparam integer d129 = 17;
        for (n129 = 0; n129 < 16; n129 = n129 + 1) 
        begin: outbit129
            assign data_11[n129 + d129*16 + c4*28*16] = data_11_array[c4][d129][n129];
        end
    endgenerate
    generate 
        localparam integer d130 = 18;
        for (n130 = 0; n130 < 16; n130 = n130 + 1) 
        begin: outbit130
            assign data_11[n130 + d130*16 + c4*28*16] = data_11_array[c4][d130][n130];
        end
    endgenerate
    generate 
        localparam integer d131 = 19;
        for (n131 = 0; n131 < 16; n131 = n131 + 1) 
        begin: outbit131
            assign data_11[n131 + d131*16 + c4*28*16] = data_11_array[c4][d131][n131];
        end
    endgenerate
    generate 
        localparam integer d132 = 20;
        for (n132 = 0; n132 < 16; n132 = n132 + 1) 
        begin: outbit132
            assign data_11[n132 + d132*16 + c4*28*16] = data_11_array[c4][d132][n132];
        end
    endgenerate
    generate 
        localparam integer d133 = 21;
        for (n133 = 0; n133 < 16; n133 = n133 + 1) 
        begin: outbit133
            assign data_11[n133 + d133*16 + c4*28*16] = data_11_array[c4][d133][n133];
        end
    endgenerate
    generate 
        localparam integer d134 = 22;
        for (n134 = 0; n134 < 16; n134 = n134 + 1) 
        begin: outbit134
            assign data_11[n134 + d134*16 + c4*28*16] = data_11_array[c4][d134][n134];
        end
    endgenerate
    generate 
        localparam integer d135 = 23;
        for (n135 = 0; n135 < 16; n135 = n135 + 1) 
        begin: outbit135
            assign data_11[n135 + d135*16 + c4*28*16] = data_11_array[c4][d135][n135];
        end
    endgenerate
    generate 
        localparam integer d136 = 24;
        for (n136 = 0; n136 < 16; n136 = n136 + 1) 
        begin: outbit136
            assign data_11[n136 + d136*16 + c4*28*16] = data_11_array[c4][d136][n136];
        end
    endgenerate
    generate 
        localparam integer d137 = 25;
        for (n137 = 0; n137 < 16; n137 = n137 + 1) 
        begin: outbit137
            assign data_11[n137 + d137*16 + c4*28*16] = data_11_array[c4][d137][n137];
        end
    endgenerate
    generate 
        localparam integer d138 = 26;
        for (n138 = 0; n138 < 16; n138 = n138 + 1) 
        begin: outbit138
            assign data_11[n138 + d138*16 + c4*28*16] = data_11_array[c4][d138][n138];
        end
    endgenerate
    generate 
        localparam integer d139 = 27;
        for (n139 = 0; n139 < 16; n139 = n139 + 1) 
        begin: outbit139
            assign data_11[n139 + d139*16 + c4*28*16] = data_11_array[c4][d139][n139];
        end
    endgenerate
    localparam integer c5 = 5;
    generate 
        localparam integer d140 = 0;
        for (n140 = 0; n140 < 16; n140 = n140 + 1) 
        begin: outbit140
            assign data_11[n140 + d140*16 + c5*28*16] = data_11_array[c5][d140][n140];
        end
    endgenerate
    generate 
        localparam integer d141 = 1;
        for (n141 = 0; n141 < 16; n141 = n141 + 1) 
        begin: outbit141
            assign data_11[n141 + d141*16 + c5*28*16] = data_11_array[c5][d141][n141];
        end
    endgenerate
    generate 
        localparam integer d142 = 2;
        for (n142 = 0; n142 < 16; n142 = n142 + 1) 
        begin: outbit142
            assign data_11[n142 + d142*16 + c5*28*16] = data_11_array[c5][d142][n142];
        end
    endgenerate
    generate 
        localparam integer d143 = 3;
        for (n143 = 0; n143 < 16; n143 = n143 + 1) 
        begin: outbit143
            assign data_11[n143 + d143*16 + c5*28*16] = data_11_array[c5][d143][n143];
        end
    endgenerate
    generate 
        localparam integer d144 = 4;
        for (n144 = 0; n144 < 16; n144 = n144 + 1) 
        begin: outbit144
            assign data_11[n144 + d144*16 + c5*28*16] = data_11_array[c5][d144][n144];
        end
    endgenerate
    generate 
        localparam integer d145 = 5;
        for (n145 = 0; n145 < 16; n145 = n145 + 1) 
        begin: outbit145
            assign data_11[n145 + d145*16 + c5*28*16] = data_11_array[c5][d145][n145];
        end
    endgenerate
    generate 
        localparam integer d146 = 6;
        for (n146 = 0; n146 < 16; n146 = n146 + 1) 
        begin: outbit146
            assign data_11[n146 + d146*16 + c5*28*16] = data_11_array[c5][d146][n146];
        end
    endgenerate
    generate 
        localparam integer d147 = 7;
        for (n147 = 0; n147 < 16; n147 = n147 + 1) 
        begin: outbit147
            assign data_11[n147 + d147*16 + c5*28*16] = data_11_array[c5][d147][n147];
        end
    endgenerate
    generate 
        localparam integer d148 = 8;
        for (n148 = 0; n148 < 16; n148 = n148 + 1) 
        begin: outbit148
            assign data_11[n148 + d148*16 + c5*28*16] = data_11_array[c5][d148][n148];
        end
    endgenerate
    generate 
        localparam integer d149 = 9;
        for (n149 = 0; n149 < 16; n149 = n149 + 1) 
        begin: outbit149
            assign data_11[n149 + d149*16 + c5*28*16] = data_11_array[c5][d149][n149];
        end
    endgenerate
    generate 
        localparam integer d150 = 10;
        for (n150 = 0; n150 < 16; n150 = n150 + 1) 
        begin: outbit150
            assign data_11[n150 + d150*16 + c5*28*16] = data_11_array[c5][d150][n150];
        end
    endgenerate
    generate 
        localparam integer d151 = 11;
        for (n151 = 0; n151 < 16; n151 = n151 + 1) 
        begin: outbit151
            assign data_11[n151 + d151*16 + c5*28*16] = data_11_array[c5][d151][n151];
        end
    endgenerate
    generate 
        localparam integer d152 = 12;
        for (n152 = 0; n152 < 16; n152 = n152 + 1) 
        begin: outbit152
            assign data_11[n152 + d152*16 + c5*28*16] = data_11_array[c5][d152][n152];
        end
    endgenerate
    generate 
        localparam integer d153 = 13;
        for (n153 = 0; n153 < 16; n153 = n153 + 1) 
        begin: outbit153
            assign data_11[n153 + d153*16 + c5*28*16] = data_11_array[c5][d153][n153];
        end
    endgenerate
    generate 
        localparam integer d154 = 14;
        for (n154 = 0; n154 < 16; n154 = n154 + 1) 
        begin: outbit154
            assign data_11[n154 + d154*16 + c5*28*16] = data_11_array[c5][d154][n154];
        end
    endgenerate
    generate 
        localparam integer d155 = 15;
        for (n155 = 0; n155 < 16; n155 = n155 + 1) 
        begin: outbit155
            assign data_11[n155 + d155*16 + c5*28*16] = data_11_array[c5][d155][n155];
        end
    endgenerate
    generate 
        localparam integer d156 = 16;
        for (n156 = 0; n156 < 16; n156 = n156 + 1) 
        begin: outbit156
            assign data_11[n156 + d156*16 + c5*28*16] = data_11_array[c5][d156][n156];
        end
    endgenerate
    generate 
        localparam integer d157 = 17;
        for (n157 = 0; n157 < 16; n157 = n157 + 1) 
        begin: outbit157
            assign data_11[n157 + d157*16 + c5*28*16] = data_11_array[c5][d157][n157];
        end
    endgenerate
    generate 
        localparam integer d158 = 18;
        for (n158 = 0; n158 < 16; n158 = n158 + 1) 
        begin: outbit158
            assign data_11[n158 + d158*16 + c5*28*16] = data_11_array[c5][d158][n158];
        end
    endgenerate
    generate 
        localparam integer d159 = 19;
        for (n159 = 0; n159 < 16; n159 = n159 + 1) 
        begin: outbit159
            assign data_11[n159 + d159*16 + c5*28*16] = data_11_array[c5][d159][n159];
        end
    endgenerate
    generate 
        localparam integer d160 = 20;
        for (n160 = 0; n160 < 16; n160 = n160 + 1) 
        begin: outbit160
            assign data_11[n160 + d160*16 + c5*28*16] = data_11_array[c5][d160][n160];
        end
    endgenerate
    generate 
        localparam integer d161 = 21;
        for (n161 = 0; n161 < 16; n161 = n161 + 1) 
        begin: outbit161
            assign data_11[n161 + d161*16 + c5*28*16] = data_11_array[c5][d161][n161];
        end
    endgenerate
    generate 
        localparam integer d162 = 22;
        for (n162 = 0; n162 < 16; n162 = n162 + 1) 
        begin: outbit162
            assign data_11[n162 + d162*16 + c5*28*16] = data_11_array[c5][d162][n162];
        end
    endgenerate
    generate 
        localparam integer d163 = 23;
        for (n163 = 0; n163 < 16; n163 = n163 + 1) 
        begin: outbit163
            assign data_11[n163 + d163*16 + c5*28*16] = data_11_array[c5][d163][n163];
        end
    endgenerate
    generate 
        localparam integer d164 = 24;
        for (n164 = 0; n164 < 16; n164 = n164 + 1) 
        begin: outbit164
            assign data_11[n164 + d164*16 + c5*28*16] = data_11_array[c5][d164][n164];
        end
    endgenerate
    generate 
        localparam integer d165 = 25;
        for (n165 = 0; n165 < 16; n165 = n165 + 1) 
        begin: outbit165
            assign data_11[n165 + d165*16 + c5*28*16] = data_11_array[c5][d165][n165];
        end
    endgenerate
    generate 
        localparam integer d166 = 26;
        for (n166 = 0; n166 < 16; n166 = n166 + 1) 
        begin: outbit166
            assign data_11[n166 + d166*16 + c5*28*16] = data_11_array[c5][d166][n166];
        end
    endgenerate
    generate 
        localparam integer d167 = 27;
        for (n167 = 0; n167 < 16; n167 = n167 + 1) 
        begin: outbit167
            assign data_11[n167 + d167*16 + c5*28*16] = data_11_array[c5][d167][n167];
        end
    endgenerate
    localparam integer c6 = 6;
    generate 
        localparam integer d168 = 0;
        for (n168 = 0; n168 < 16; n168 = n168 + 1) 
        begin: outbit168
            assign data_11[n168 + d168*16 + c6*28*16] = data_11_array[c6][d168][n168];
        end
    endgenerate
    generate 
        localparam integer d169 = 1;
        for (n169 = 0; n169 < 16; n169 = n169 + 1) 
        begin: outbit169
            assign data_11[n169 + d169*16 + c6*28*16] = data_11_array[c6][d169][n169];
        end
    endgenerate
    generate 
        localparam integer d170 = 2;
        for (n170 = 0; n170 < 16; n170 = n170 + 1) 
        begin: outbit170
            assign data_11[n170 + d170*16 + c6*28*16] = data_11_array[c6][d170][n170];
        end
    endgenerate
    generate 
        localparam integer d171 = 3;
        for (n171 = 0; n171 < 16; n171 = n171 + 1) 
        begin: outbit171
            assign data_11[n171 + d171*16 + c6*28*16] = data_11_array[c6][d171][n171];
        end
    endgenerate
    generate 
        localparam integer d172 = 4;
        for (n172 = 0; n172 < 16; n172 = n172 + 1) 
        begin: outbit172
            assign data_11[n172 + d172*16 + c6*28*16] = data_11_array[c6][d172][n172];
        end
    endgenerate
    generate 
        localparam integer d173 = 5;
        for (n173 = 0; n173 < 16; n173 = n173 + 1) 
        begin: outbit173
            assign data_11[n173 + d173*16 + c6*28*16] = data_11_array[c6][d173][n173];
        end
    endgenerate
    generate 
        localparam integer d174 = 6;
        for (n174 = 0; n174 < 16; n174 = n174 + 1) 
        begin: outbit174
            assign data_11[n174 + d174*16 + c6*28*16] = data_11_array[c6][d174][n174];
        end
    endgenerate
    generate 
        localparam integer d175 = 7;
        for (n175 = 0; n175 < 16; n175 = n175 + 1) 
        begin: outbit175
            assign data_11[n175 + d175*16 + c6*28*16] = data_11_array[c6][d175][n175];
        end
    endgenerate
    generate 
        localparam integer d176 = 8;
        for (n176 = 0; n176 < 16; n176 = n176 + 1) 
        begin: outbit176
            assign data_11[n176 + d176*16 + c6*28*16] = data_11_array[c6][d176][n176];
        end
    endgenerate
    generate 
        localparam integer d177 = 9;
        for (n177 = 0; n177 < 16; n177 = n177 + 1) 
        begin: outbit177
            assign data_11[n177 + d177*16 + c6*28*16] = data_11_array[c6][d177][n177];
        end
    endgenerate
    generate 
        localparam integer d178 = 10;
        for (n178 = 0; n178 < 16; n178 = n178 + 1) 
        begin: outbit178
            assign data_11[n178 + d178*16 + c6*28*16] = data_11_array[c6][d178][n178];
        end
    endgenerate
    generate 
        localparam integer d179 = 11;
        for (n179 = 0; n179 < 16; n179 = n179 + 1) 
        begin: outbit179
            assign data_11[n179 + d179*16 + c6*28*16] = data_11_array[c6][d179][n179];
        end
    endgenerate
    generate 
        localparam integer d180 = 12;
        for (n180 = 0; n180 < 16; n180 = n180 + 1) 
        begin: outbit180
            assign data_11[n180 + d180*16 + c6*28*16] = data_11_array[c6][d180][n180];
        end
    endgenerate
    generate 
        localparam integer d181 = 13;
        for (n181 = 0; n181 < 16; n181 = n181 + 1) 
        begin: outbit181
            assign data_11[n181 + d181*16 + c6*28*16] = data_11_array[c6][d181][n181];
        end
    endgenerate
    generate 
        localparam integer d182 = 14;
        for (n182 = 0; n182 < 16; n182 = n182 + 1) 
        begin: outbit182
            assign data_11[n182 + d182*16 + c6*28*16] = data_11_array[c6][d182][n182];
        end
    endgenerate
    generate 
        localparam integer d183 = 15;
        for (n183 = 0; n183 < 16; n183 = n183 + 1) 
        begin: outbit183
            assign data_11[n183 + d183*16 + c6*28*16] = data_11_array[c6][d183][n183];
        end
    endgenerate
    generate 
        localparam integer d184 = 16;
        for (n184 = 0; n184 < 16; n184 = n184 + 1) 
        begin: outbit184
            assign data_11[n184 + d184*16 + c6*28*16] = data_11_array[c6][d184][n184];
        end
    endgenerate
    generate 
        localparam integer d185 = 17;
        for (n185 = 0; n185 < 16; n185 = n185 + 1) 
        begin: outbit185
            assign data_11[n185 + d185*16 + c6*28*16] = data_11_array[c6][d185][n185];
        end
    endgenerate
    generate 
        localparam integer d186 = 18;
        for (n186 = 0; n186 < 16; n186 = n186 + 1) 
        begin: outbit186
            assign data_11[n186 + d186*16 + c6*28*16] = data_11_array[c6][d186][n186];
        end
    endgenerate
    generate 
        localparam integer d187 = 19;
        for (n187 = 0; n187 < 16; n187 = n187 + 1) 
        begin: outbit187
            assign data_11[n187 + d187*16 + c6*28*16] = data_11_array[c6][d187][n187];
        end
    endgenerate
    generate 
        localparam integer d188 = 20;
        for (n188 = 0; n188 < 16; n188 = n188 + 1) 
        begin: outbit188
            assign data_11[n188 + d188*16 + c6*28*16] = data_11_array[c6][d188][n188];
        end
    endgenerate
    generate 
        localparam integer d189 = 21;
        for (n189 = 0; n189 < 16; n189 = n189 + 1) 
        begin: outbit189
            assign data_11[n189 + d189*16 + c6*28*16] = data_11_array[c6][d189][n189];
        end
    endgenerate
    generate 
        localparam integer d190 = 22;
        for (n190 = 0; n190 < 16; n190 = n190 + 1) 
        begin: outbit190
            assign data_11[n190 + d190*16 + c6*28*16] = data_11_array[c6][d190][n190];
        end
    endgenerate
    generate 
        localparam integer d191 = 23;
        for (n191 = 0; n191 < 16; n191 = n191 + 1) 
        begin: outbit191
            assign data_11[n191 + d191*16 + c6*28*16] = data_11_array[c6][d191][n191];
        end
    endgenerate
    generate 
        localparam integer d192 = 24;
        for (n192 = 0; n192 < 16; n192 = n192 + 1) 
        begin: outbit192
            assign data_11[n192 + d192*16 + c6*28*16] = data_11_array[c6][d192][n192];
        end
    endgenerate
    generate 
        localparam integer d193 = 25;
        for (n193 = 0; n193 < 16; n193 = n193 + 1) 
        begin: outbit193
            assign data_11[n193 + d193*16 + c6*28*16] = data_11_array[c6][d193][n193];
        end
    endgenerate
    generate 
        localparam integer d194 = 26;
        for (n194 = 0; n194 < 16; n194 = n194 + 1) 
        begin: outbit194
            assign data_11[n194 + d194*16 + c6*28*16] = data_11_array[c6][d194][n194];
        end
    endgenerate
    generate 
        localparam integer d195 = 27;
        for (n195 = 0; n195 < 16; n195 = n195 + 1) 
        begin: outbit195
            assign data_11[n195 + d195*16 + c6*28*16] = data_11_array[c6][d195][n195];
        end
    endgenerate
    localparam integer c7 = 7;
    generate 
        localparam integer d196 = 0;
        for (n196 = 0; n196 < 16; n196 = n196 + 1) 
        begin: outbit196
            assign data_11[n196 + d196*16 + c7*28*16] = data_11_array[c7][d196][n196];
        end
    endgenerate
    generate 
        localparam integer d197 = 1;
        for (n197 = 0; n197 < 16; n197 = n197 + 1) 
        begin: outbit197
            assign data_11[n197 + d197*16 + c7*28*16] = data_11_array[c7][d197][n197];
        end
    endgenerate
    generate 
        localparam integer d198 = 2;
        for (n198 = 0; n198 < 16; n198 = n198 + 1) 
        begin: outbit198
            assign data_11[n198 + d198*16 + c7*28*16] = data_11_array[c7][d198][n198];
        end
    endgenerate
    generate 
        localparam integer d199 = 3;
        for (n199 = 0; n199 < 16; n199 = n199 + 1) 
        begin: outbit199
            assign data_11[n199 + d199*16 + c7*28*16] = data_11_array[c7][d199][n199];
        end
    endgenerate
    generate 
        localparam integer d200 = 4;
        for (n200 = 0; n200 < 16; n200 = n200 + 1) 
        begin: outbit200
            assign data_11[n200 + d200*16 + c7*28*16] = data_11_array[c7][d200][n200];
        end
    endgenerate
    generate 
        localparam integer d201 = 5;
        for (n201 = 0; n201 < 16; n201 = n201 + 1) 
        begin: outbit201
            assign data_11[n201 + d201*16 + c7*28*16] = data_11_array[c7][d201][n201];
        end
    endgenerate
    generate 
        localparam integer d202 = 6;
        for (n202 = 0; n202 < 16; n202 = n202 + 1) 
        begin: outbit202
            assign data_11[n202 + d202*16 + c7*28*16] = data_11_array[c7][d202][n202];
        end
    endgenerate
    generate 
        localparam integer d203 = 7;
        for (n203 = 0; n203 < 16; n203 = n203 + 1) 
        begin: outbit203
            assign data_11[n203 + d203*16 + c7*28*16] = data_11_array[c7][d203][n203];
        end
    endgenerate
    generate 
        localparam integer d204 = 8;
        for (n204 = 0; n204 < 16; n204 = n204 + 1) 
        begin: outbit204
            assign data_11[n204 + d204*16 + c7*28*16] = data_11_array[c7][d204][n204];
        end
    endgenerate
    generate 
        localparam integer d205 = 9;
        for (n205 = 0; n205 < 16; n205 = n205 + 1) 
        begin: outbit205
            assign data_11[n205 + d205*16 + c7*28*16] = data_11_array[c7][d205][n205];
        end
    endgenerate
    generate 
        localparam integer d206 = 10;
        for (n206 = 0; n206 < 16; n206 = n206 + 1) 
        begin: outbit206
            assign data_11[n206 + d206*16 + c7*28*16] = data_11_array[c7][d206][n206];
        end
    endgenerate
    generate 
        localparam integer d207 = 11;
        for (n207 = 0; n207 < 16; n207 = n207 + 1) 
        begin: outbit207
            assign data_11[n207 + d207*16 + c7*28*16] = data_11_array[c7][d207][n207];
        end
    endgenerate
    generate 
        localparam integer d208 = 12;
        for (n208 = 0; n208 < 16; n208 = n208 + 1) 
        begin: outbit208
            assign data_11[n208 + d208*16 + c7*28*16] = data_11_array[c7][d208][n208];
        end
    endgenerate
    generate 
        localparam integer d209 = 13;
        for (n209 = 0; n209 < 16; n209 = n209 + 1) 
        begin: outbit209
            assign data_11[n209 + d209*16 + c7*28*16] = data_11_array[c7][d209][n209];
        end
    endgenerate
    generate 
        localparam integer d210 = 14;
        for (n210 = 0; n210 < 16; n210 = n210 + 1) 
        begin: outbit210
            assign data_11[n210 + d210*16 + c7*28*16] = data_11_array[c7][d210][n210];
        end
    endgenerate
    generate 
        localparam integer d211 = 15;
        for (n211 = 0; n211 < 16; n211 = n211 + 1) 
        begin: outbit211
            assign data_11[n211 + d211*16 + c7*28*16] = data_11_array[c7][d211][n211];
        end
    endgenerate
    generate 
        localparam integer d212 = 16;
        for (n212 = 0; n212 < 16; n212 = n212 + 1) 
        begin: outbit212
            assign data_11[n212 + d212*16 + c7*28*16] = data_11_array[c7][d212][n212];
        end
    endgenerate
    generate 
        localparam integer d213 = 17;
        for (n213 = 0; n213 < 16; n213 = n213 + 1) 
        begin: outbit213
            assign data_11[n213 + d213*16 + c7*28*16] = data_11_array[c7][d213][n213];
        end
    endgenerate
    generate 
        localparam integer d214 = 18;
        for (n214 = 0; n214 < 16; n214 = n214 + 1) 
        begin: outbit214
            assign data_11[n214 + d214*16 + c7*28*16] = data_11_array[c7][d214][n214];
        end
    endgenerate
    generate 
        localparam integer d215 = 19;
        for (n215 = 0; n215 < 16; n215 = n215 + 1) 
        begin: outbit215
            assign data_11[n215 + d215*16 + c7*28*16] = data_11_array[c7][d215][n215];
        end
    endgenerate
    generate 
        localparam integer d216 = 20;
        for (n216 = 0; n216 < 16; n216 = n216 + 1) 
        begin: outbit216
            assign data_11[n216 + d216*16 + c7*28*16] = data_11_array[c7][d216][n216];
        end
    endgenerate
    generate 
        localparam integer d217 = 21;
        for (n217 = 0; n217 < 16; n217 = n217 + 1) 
        begin: outbit217
            assign data_11[n217 + d217*16 + c7*28*16] = data_11_array[c7][d217][n217];
        end
    endgenerate
    generate 
        localparam integer d218 = 22;
        for (n218 = 0; n218 < 16; n218 = n218 + 1) 
        begin: outbit218
            assign data_11[n218 + d218*16 + c7*28*16] = data_11_array[c7][d218][n218];
        end
    endgenerate
    generate 
        localparam integer d219 = 23;
        for (n219 = 0; n219 < 16; n219 = n219 + 1) 
        begin: outbit219
            assign data_11[n219 + d219*16 + c7*28*16] = data_11_array[c7][d219][n219];
        end
    endgenerate
    generate 
        localparam integer d220 = 24;
        for (n220 = 0; n220 < 16; n220 = n220 + 1) 
        begin: outbit220
            assign data_11[n220 + d220*16 + c7*28*16] = data_11_array[c7][d220][n220];
        end
    endgenerate
    generate 
        localparam integer d221 = 25;
        for (n221 = 0; n221 < 16; n221 = n221 + 1) 
        begin: outbit221
            assign data_11[n221 + d221*16 + c7*28*16] = data_11_array[c7][d221][n221];
        end
    endgenerate
    generate 
        localparam integer d222 = 26;
        for (n222 = 0; n222 < 16; n222 = n222 + 1) 
        begin: outbit222
            assign data_11[n222 + d222*16 + c7*28*16] = data_11_array[c7][d222][n222];
        end
    endgenerate
    generate 
        localparam integer d223 = 27;
        for (n223 = 0; n223 < 16; n223 = n223 + 1) 
        begin: outbit223
            assign data_11[n223 + d223*16 + c7*28*16] = data_11_array[c7][d223][n223];
        end
    endgenerate
    localparam integer c8 = 8;
    generate 
        localparam integer d224 = 0;
        for (n224 = 0; n224 < 16; n224 = n224 + 1) 
        begin: outbit224
            assign data_11[n224 + d224*16 + c8*28*16] = data_11_array[c8][d224][n224];
        end
    endgenerate
    generate 
        localparam integer d225 = 1;
        for (n225 = 0; n225 < 16; n225 = n225 + 1) 
        begin: outbit225
            assign data_11[n225 + d225*16 + c8*28*16] = data_11_array[c8][d225][n225];
        end
    endgenerate
    generate 
        localparam integer d226 = 2;
        for (n226 = 0; n226 < 16; n226 = n226 + 1) 
        begin: outbit226
            assign data_11[n226 + d226*16 + c8*28*16] = data_11_array[c8][d226][n226];
        end
    endgenerate
    generate 
        localparam integer d227 = 3;
        for (n227 = 0; n227 < 16; n227 = n227 + 1) 
        begin: outbit227
            assign data_11[n227 + d227*16 + c8*28*16] = data_11_array[c8][d227][n227];
        end
    endgenerate
    generate 
        localparam integer d228 = 4;
        for (n228 = 0; n228 < 16; n228 = n228 + 1) 
        begin: outbit228
            assign data_11[n228 + d228*16 + c8*28*16] = data_11_array[c8][d228][n228];
        end
    endgenerate
    generate 
        localparam integer d229 = 5;
        for (n229 = 0; n229 < 16; n229 = n229 + 1) 
        begin: outbit229
            assign data_11[n229 + d229*16 + c8*28*16] = data_11_array[c8][d229][n229];
        end
    endgenerate
    generate 
        localparam integer d230 = 6;
        for (n230 = 0; n230 < 16; n230 = n230 + 1) 
        begin: outbit230
            assign data_11[n230 + d230*16 + c8*28*16] = data_11_array[c8][d230][n230];
        end
    endgenerate
    generate 
        localparam integer d231 = 7;
        for (n231 = 0; n231 < 16; n231 = n231 + 1) 
        begin: outbit231
            assign data_11[n231 + d231*16 + c8*28*16] = data_11_array[c8][d231][n231];
        end
    endgenerate
    generate 
        localparam integer d232 = 8;
        for (n232 = 0; n232 < 16; n232 = n232 + 1) 
        begin: outbit232
            assign data_11[n232 + d232*16 + c8*28*16] = data_11_array[c8][d232][n232];
        end
    endgenerate
    generate 
        localparam integer d233 = 9;
        for (n233 = 0; n233 < 16; n233 = n233 + 1) 
        begin: outbit233
            assign data_11[n233 + d233*16 + c8*28*16] = data_11_array[c8][d233][n233];
        end
    endgenerate
    generate 
        localparam integer d234 = 10;
        for (n234 = 0; n234 < 16; n234 = n234 + 1) 
        begin: outbit234
            assign data_11[n234 + d234*16 + c8*28*16] = data_11_array[c8][d234][n234];
        end
    endgenerate
    generate 
        localparam integer d235 = 11;
        for (n235 = 0; n235 < 16; n235 = n235 + 1) 
        begin: outbit235
            assign data_11[n235 + d235*16 + c8*28*16] = data_11_array[c8][d235][n235];
        end
    endgenerate
    generate 
        localparam integer d236 = 12;
        for (n236 = 0; n236 < 16; n236 = n236 + 1) 
        begin: outbit236
            assign data_11[n236 + d236*16 + c8*28*16] = data_11_array[c8][d236][n236];
        end
    endgenerate
    generate 
        localparam integer d237 = 13;
        for (n237 = 0; n237 < 16; n237 = n237 + 1) 
        begin: outbit237
            assign data_11[n237 + d237*16 + c8*28*16] = data_11_array[c8][d237][n237];
        end
    endgenerate
    generate 
        localparam integer d238 = 14;
        for (n238 = 0; n238 < 16; n238 = n238 + 1) 
        begin: outbit238
            assign data_11[n238 + d238*16 + c8*28*16] = data_11_array[c8][d238][n238];
        end
    endgenerate
    generate 
        localparam integer d239 = 15;
        for (n239 = 0; n239 < 16; n239 = n239 + 1) 
        begin: outbit239
            assign data_11[n239 + d239*16 + c8*28*16] = data_11_array[c8][d239][n239];
        end
    endgenerate
    generate 
        localparam integer d240 = 16;
        for (n240 = 0; n240 < 16; n240 = n240 + 1) 
        begin: outbit240
            assign data_11[n240 + d240*16 + c8*28*16] = data_11_array[c8][d240][n240];
        end
    endgenerate
    generate 
        localparam integer d241 = 17;
        for (n241 = 0; n241 < 16; n241 = n241 + 1) 
        begin: outbit241
            assign data_11[n241 + d241*16 + c8*28*16] = data_11_array[c8][d241][n241];
        end
    endgenerate
    generate 
        localparam integer d242 = 18;
        for (n242 = 0; n242 < 16; n242 = n242 + 1) 
        begin: outbit242
            assign data_11[n242 + d242*16 + c8*28*16] = data_11_array[c8][d242][n242];
        end
    endgenerate
    generate 
        localparam integer d243 = 19;
        for (n243 = 0; n243 < 16; n243 = n243 + 1) 
        begin: outbit243
            assign data_11[n243 + d243*16 + c8*28*16] = data_11_array[c8][d243][n243];
        end
    endgenerate
    generate 
        localparam integer d244 = 20;
        for (n244 = 0; n244 < 16; n244 = n244 + 1) 
        begin: outbit244
            assign data_11[n244 + d244*16 + c8*28*16] = data_11_array[c8][d244][n244];
        end
    endgenerate
    generate 
        localparam integer d245 = 21;
        for (n245 = 0; n245 < 16; n245 = n245 + 1) 
        begin: outbit245
            assign data_11[n245 + d245*16 + c8*28*16] = data_11_array[c8][d245][n245];
        end
    endgenerate
    generate 
        localparam integer d246 = 22;
        for (n246 = 0; n246 < 16; n246 = n246 + 1) 
        begin: outbit246
            assign data_11[n246 + d246*16 + c8*28*16] = data_11_array[c8][d246][n246];
        end
    endgenerate
    generate 
        localparam integer d247 = 23;
        for (n247 = 0; n247 < 16; n247 = n247 + 1) 
        begin: outbit247
            assign data_11[n247 + d247*16 + c8*28*16] = data_11_array[c8][d247][n247];
        end
    endgenerate
    generate 
        localparam integer d248 = 24;
        for (n248 = 0; n248 < 16; n248 = n248 + 1) 
        begin: outbit248
            assign data_11[n248 + d248*16 + c8*28*16] = data_11_array[c8][d248][n248];
        end
    endgenerate
    generate 
        localparam integer d249 = 25;
        for (n249 = 0; n249 < 16; n249 = n249 + 1) 
        begin: outbit249
            assign data_11[n249 + d249*16 + c8*28*16] = data_11_array[c8][d249][n249];
        end
    endgenerate
    generate 
        localparam integer d250 = 26;
        for (n250 = 0; n250 < 16; n250 = n250 + 1) 
        begin: outbit250
            assign data_11[n250 + d250*16 + c8*28*16] = data_11_array[c8][d250][n250];
        end
    endgenerate
    generate 
        localparam integer d251 = 27;
        for (n251 = 0; n251 < 16; n251 = n251 + 1) 
        begin: outbit251
            assign data_11[n251 + d251*16 + c8*28*16] = data_11_array[c8][d251][n251];
        end
    endgenerate
    localparam integer c9 = 9;
    generate 
        localparam integer d252 = 0;
        for (n252 = 0; n252 < 16; n252 = n252 + 1) 
        begin: outbit252
            assign data_11[n252 + d252*16 + c9*28*16] = data_11_array[c9][d252][n252];
        end
    endgenerate
    generate 
        localparam integer d253 = 1;
        for (n253 = 0; n253 < 16; n253 = n253 + 1) 
        begin: outbit253
            assign data_11[n253 + d253*16 + c9*28*16] = data_11_array[c9][d253][n253];
        end
    endgenerate
    generate 
        localparam integer d254 = 2;
        for (n254 = 0; n254 < 16; n254 = n254 + 1) 
        begin: outbit254
            assign data_11[n254 + d254*16 + c9*28*16] = data_11_array[c9][d254][n254];
        end
    endgenerate
    generate 
        localparam integer d255 = 3;
        for (n255 = 0; n255 < 16; n255 = n255 + 1) 
        begin: outbit255
            assign data_11[n255 + d255*16 + c9*28*16] = data_11_array[c9][d255][n255];
        end
    endgenerate
    generate 
        localparam integer d256 = 4;
        for (n256 = 0; n256 < 16; n256 = n256 + 1) 
        begin: outbit256
            assign data_11[n256 + d256*16 + c9*28*16] = data_11_array[c9][d256][n256];
        end
    endgenerate
    generate 
        localparam integer d257 = 5;
        for (n257 = 0; n257 < 16; n257 = n257 + 1) 
        begin: outbit257
            assign data_11[n257 + d257*16 + c9*28*16] = data_11_array[c9][d257][n257];
        end
    endgenerate
    generate 
        localparam integer d258 = 6;
        for (n258 = 0; n258 < 16; n258 = n258 + 1) 
        begin: outbit258
            assign data_11[n258 + d258*16 + c9*28*16] = data_11_array[c9][d258][n258];
        end
    endgenerate
    generate 
        localparam integer d259 = 7;
        for (n259 = 0; n259 < 16; n259 = n259 + 1) 
        begin: outbit259
            assign data_11[n259 + d259*16 + c9*28*16] = data_11_array[c9][d259][n259];
        end
    endgenerate
    generate 
        localparam integer d260 = 8;
        for (n260 = 0; n260 < 16; n260 = n260 + 1) 
        begin: outbit260
            assign data_11[n260 + d260*16 + c9*28*16] = data_11_array[c9][d260][n260];
        end
    endgenerate
    generate 
        localparam integer d261 = 9;
        for (n261 = 0; n261 < 16; n261 = n261 + 1) 
        begin: outbit261
            assign data_11[n261 + d261*16 + c9*28*16] = data_11_array[c9][d261][n261];
        end
    endgenerate
    generate 
        localparam integer d262 = 10;
        for (n262 = 0; n262 < 16; n262 = n262 + 1) 
        begin: outbit262
            assign data_11[n262 + d262*16 + c9*28*16] = data_11_array[c9][d262][n262];
        end
    endgenerate
    generate 
        localparam integer d263 = 11;
        for (n263 = 0; n263 < 16; n263 = n263 + 1) 
        begin: outbit263
            assign data_11[n263 + d263*16 + c9*28*16] = data_11_array[c9][d263][n263];
        end
    endgenerate
    generate 
        localparam integer d264 = 12;
        for (n264 = 0; n264 < 16; n264 = n264 + 1) 
        begin: outbit264
            assign data_11[n264 + d264*16 + c9*28*16] = data_11_array[c9][d264][n264];
        end
    endgenerate
    generate 
        localparam integer d265 = 13;
        for (n265 = 0; n265 < 16; n265 = n265 + 1) 
        begin: outbit265
            assign data_11[n265 + d265*16 + c9*28*16] = data_11_array[c9][d265][n265];
        end
    endgenerate
    generate 
        localparam integer d266 = 14;
        for (n266 = 0; n266 < 16; n266 = n266 + 1) 
        begin: outbit266
            assign data_11[n266 + d266*16 + c9*28*16] = data_11_array[c9][d266][n266];
        end
    endgenerate
    generate 
        localparam integer d267 = 15;
        for (n267 = 0; n267 < 16; n267 = n267 + 1) 
        begin: outbit267
            assign data_11[n267 + d267*16 + c9*28*16] = data_11_array[c9][d267][n267];
        end
    endgenerate
    generate 
        localparam integer d268 = 16;
        for (n268 = 0; n268 < 16; n268 = n268 + 1) 
        begin: outbit268
            assign data_11[n268 + d268*16 + c9*28*16] = data_11_array[c9][d268][n268];
        end
    endgenerate
    generate 
        localparam integer d269 = 17;
        for (n269 = 0; n269 < 16; n269 = n269 + 1) 
        begin: outbit269
            assign data_11[n269 + d269*16 + c9*28*16] = data_11_array[c9][d269][n269];
        end
    endgenerate
    generate 
        localparam integer d270 = 18;
        for (n270 = 0; n270 < 16; n270 = n270 + 1) 
        begin: outbit270
            assign data_11[n270 + d270*16 + c9*28*16] = data_11_array[c9][d270][n270];
        end
    endgenerate
    generate 
        localparam integer d271 = 19;
        for (n271 = 0; n271 < 16; n271 = n271 + 1) 
        begin: outbit271
            assign data_11[n271 + d271*16 + c9*28*16] = data_11_array[c9][d271][n271];
        end
    endgenerate
    generate 
        localparam integer d272 = 20;
        for (n272 = 0; n272 < 16; n272 = n272 + 1) 
        begin: outbit272
            assign data_11[n272 + d272*16 + c9*28*16] = data_11_array[c9][d272][n272];
        end
    endgenerate
    generate 
        localparam integer d273 = 21;
        for (n273 = 0; n273 < 16; n273 = n273 + 1) 
        begin: outbit273
            assign data_11[n273 + d273*16 + c9*28*16] = data_11_array[c9][d273][n273];
        end
    endgenerate
    generate 
        localparam integer d274 = 22;
        for (n274 = 0; n274 < 16; n274 = n274 + 1) 
        begin: outbit274
            assign data_11[n274 + d274*16 + c9*28*16] = data_11_array[c9][d274][n274];
        end
    endgenerate
    generate 
        localparam integer d275 = 23;
        for (n275 = 0; n275 < 16; n275 = n275 + 1) 
        begin: outbit275
            assign data_11[n275 + d275*16 + c9*28*16] = data_11_array[c9][d275][n275];
        end
    endgenerate
    generate 
        localparam integer d276 = 24;
        for (n276 = 0; n276 < 16; n276 = n276 + 1) 
        begin: outbit276
            assign data_11[n276 + d276*16 + c9*28*16] = data_11_array[c9][d276][n276];
        end
    endgenerate
    generate 
        localparam integer d277 = 25;
        for (n277 = 0; n277 < 16; n277 = n277 + 1) 
        begin: outbit277
            assign data_11[n277 + d277*16 + c9*28*16] = data_11_array[c9][d277][n277];
        end
    endgenerate
    generate 
        localparam integer d278 = 26;
        for (n278 = 0; n278 < 16; n278 = n278 + 1) 
        begin: outbit278
            assign data_11[n278 + d278*16 + c9*28*16] = data_11_array[c9][d278][n278];
        end
    endgenerate
    generate 
        localparam integer d279 = 27;
        for (n279 = 0; n279 < 16; n279 = n279 + 1) 
        begin: outbit279
            assign data_11[n279 + d279*16 + c9*28*16] = data_11_array[c9][d279][n279];
        end
    endgenerate
    localparam integer c10 = 10;
    generate 
        localparam integer d280 = 0;
        for (n280 = 0; n280 < 16; n280 = n280 + 1) 
        begin: outbit280
            assign data_11[n280 + d280*16 + c10*28*16] = data_11_array[c10][d280][n280];
        end
    endgenerate
    generate 
        localparam integer d281 = 1;
        for (n281 = 0; n281 < 16; n281 = n281 + 1) 
        begin: outbit281
            assign data_11[n281 + d281*16 + c10*28*16] = data_11_array[c10][d281][n281];
        end
    endgenerate
    generate 
        localparam integer d282 = 2;
        for (n282 = 0; n282 < 16; n282 = n282 + 1) 
        begin: outbit282
            assign data_11[n282 + d282*16 + c10*28*16] = data_11_array[c10][d282][n282];
        end
    endgenerate
    generate 
        localparam integer d283 = 3;
        for (n283 = 0; n283 < 16; n283 = n283 + 1) 
        begin: outbit283
            assign data_11[n283 + d283*16 + c10*28*16] = data_11_array[c10][d283][n283];
        end
    endgenerate
    generate 
        localparam integer d284 = 4;
        for (n284 = 0; n284 < 16; n284 = n284 + 1) 
        begin: outbit284
            assign data_11[n284 + d284*16 + c10*28*16] = data_11_array[c10][d284][n284];
        end
    endgenerate
    generate 
        localparam integer d285 = 5;
        for (n285 = 0; n285 < 16; n285 = n285 + 1) 
        begin: outbit285
            assign data_11[n285 + d285*16 + c10*28*16] = data_11_array[c10][d285][n285];
        end
    endgenerate
    generate 
        localparam integer d286 = 6;
        for (n286 = 0; n286 < 16; n286 = n286 + 1) 
        begin: outbit286
            assign data_11[n286 + d286*16 + c10*28*16] = data_11_array[c10][d286][n286];
        end
    endgenerate
    generate 
        localparam integer d287 = 7;
        for (n287 = 0; n287 < 16; n287 = n287 + 1) 
        begin: outbit287
            assign data_11[n287 + d287*16 + c10*28*16] = data_11_array[c10][d287][n287];
        end
    endgenerate
    generate 
        localparam integer d288 = 8;
        for (n288 = 0; n288 < 16; n288 = n288 + 1) 
        begin: outbit288
            assign data_11[n288 + d288*16 + c10*28*16] = data_11_array[c10][d288][n288];
        end
    endgenerate
    generate 
        localparam integer d289 = 9;
        for (n289 = 0; n289 < 16; n289 = n289 + 1) 
        begin: outbit289
            assign data_11[n289 + d289*16 + c10*28*16] = data_11_array[c10][d289][n289];
        end
    endgenerate
    generate 
        localparam integer d290 = 10;
        for (n290 = 0; n290 < 16; n290 = n290 + 1) 
        begin: outbit290
            assign data_11[n290 + d290*16 + c10*28*16] = data_11_array[c10][d290][n290];
        end
    endgenerate
    generate 
        localparam integer d291 = 11;
        for (n291 = 0; n291 < 16; n291 = n291 + 1) 
        begin: outbit291
            assign data_11[n291 + d291*16 + c10*28*16] = data_11_array[c10][d291][n291];
        end
    endgenerate
    generate 
        localparam integer d292 = 12;
        for (n292 = 0; n292 < 16; n292 = n292 + 1) 
        begin: outbit292
            assign data_11[n292 + d292*16 + c10*28*16] = data_11_array[c10][d292][n292];
        end
    endgenerate
    generate 
        localparam integer d293 = 13;
        for (n293 = 0; n293 < 16; n293 = n293 + 1) 
        begin: outbit293
            assign data_11[n293 + d293*16 + c10*28*16] = data_11_array[c10][d293][n293];
        end
    endgenerate
    generate 
        localparam integer d294 = 14;
        for (n294 = 0; n294 < 16; n294 = n294 + 1) 
        begin: outbit294
            assign data_11[n294 + d294*16 + c10*28*16] = data_11_array[c10][d294][n294];
        end
    endgenerate
    generate 
        localparam integer d295 = 15;
        for (n295 = 0; n295 < 16; n295 = n295 + 1) 
        begin: outbit295
            assign data_11[n295 + d295*16 + c10*28*16] = data_11_array[c10][d295][n295];
        end
    endgenerate
    generate 
        localparam integer d296 = 16;
        for (n296 = 0; n296 < 16; n296 = n296 + 1) 
        begin: outbit296
            assign data_11[n296 + d296*16 + c10*28*16] = data_11_array[c10][d296][n296];
        end
    endgenerate
    generate 
        localparam integer d297 = 17;
        for (n297 = 0; n297 < 16; n297 = n297 + 1) 
        begin: outbit297
            assign data_11[n297 + d297*16 + c10*28*16] = data_11_array[c10][d297][n297];
        end
    endgenerate
    generate 
        localparam integer d298 = 18;
        for (n298 = 0; n298 < 16; n298 = n298 + 1) 
        begin: outbit298
            assign data_11[n298 + d298*16 + c10*28*16] = data_11_array[c10][d298][n298];
        end
    endgenerate
    generate 
        localparam integer d299 = 19;
        for (n299 = 0; n299 < 16; n299 = n299 + 1) 
        begin: outbit299
            assign data_11[n299 + d299*16 + c10*28*16] = data_11_array[c10][d299][n299];
        end
    endgenerate
    generate 
        localparam integer d300 = 20;
        for (n300 = 0; n300 < 16; n300 = n300 + 1) 
        begin: outbit300
            assign data_11[n300 + d300*16 + c10*28*16] = data_11_array[c10][d300][n300];
        end
    endgenerate
    generate 
        localparam integer d301 = 21;
        for (n301 = 0; n301 < 16; n301 = n301 + 1) 
        begin: outbit301
            assign data_11[n301 + d301*16 + c10*28*16] = data_11_array[c10][d301][n301];
        end
    endgenerate
    generate 
        localparam integer d302 = 22;
        for (n302 = 0; n302 < 16; n302 = n302 + 1) 
        begin: outbit302
            assign data_11[n302 + d302*16 + c10*28*16] = data_11_array[c10][d302][n302];
        end
    endgenerate
    generate 
        localparam integer d303 = 23;
        for (n303 = 0; n303 < 16; n303 = n303 + 1) 
        begin: outbit303
            assign data_11[n303 + d303*16 + c10*28*16] = data_11_array[c10][d303][n303];
        end
    endgenerate
    generate 
        localparam integer d304 = 24;
        for (n304 = 0; n304 < 16; n304 = n304 + 1) 
        begin: outbit304
            assign data_11[n304 + d304*16 + c10*28*16] = data_11_array[c10][d304][n304];
        end
    endgenerate
    generate 
        localparam integer d305 = 25;
        for (n305 = 0; n305 < 16; n305 = n305 + 1) 
        begin: outbit305
            assign data_11[n305 + d305*16 + c10*28*16] = data_11_array[c10][d305][n305];
        end
    endgenerate
    generate 
        localparam integer d306 = 26;
        for (n306 = 0; n306 < 16; n306 = n306 + 1) 
        begin: outbit306
            assign data_11[n306 + d306*16 + c10*28*16] = data_11_array[c10][d306][n306];
        end
    endgenerate
    generate 
        localparam integer d307 = 27;
        for (n307 = 0; n307 < 16; n307 = n307 + 1) 
        begin: outbit307
            assign data_11[n307 + d307*16 + c10*28*16] = data_11_array[c10][d307][n307];
        end
    endgenerate
    localparam integer c11 = 11;
    generate 
        localparam integer d308 = 0;
        for (n308 = 0; n308 < 16; n308 = n308 + 1) 
        begin: outbit308
            assign data_11[n308 + d308*16 + c11*28*16] = data_11_array[c11][d308][n308];
        end
    endgenerate
    generate 
        localparam integer d309 = 1;
        for (n309 = 0; n309 < 16; n309 = n309 + 1) 
        begin: outbit309
            assign data_11[n309 + d309*16 + c11*28*16] = data_11_array[c11][d309][n309];
        end
    endgenerate
    generate 
        localparam integer d310 = 2;
        for (n310 = 0; n310 < 16; n310 = n310 + 1) 
        begin: outbit310
            assign data_11[n310 + d310*16 + c11*28*16] = data_11_array[c11][d310][n310];
        end
    endgenerate
    generate 
        localparam integer d311 = 3;
        for (n311 = 0; n311 < 16; n311 = n311 + 1) 
        begin: outbit311
            assign data_11[n311 + d311*16 + c11*28*16] = data_11_array[c11][d311][n311];
        end
    endgenerate
    generate 
        localparam integer d312 = 4;
        for (n312 = 0; n312 < 16; n312 = n312 + 1) 
        begin: outbit312
            assign data_11[n312 + d312*16 + c11*28*16] = data_11_array[c11][d312][n312];
        end
    endgenerate
    generate 
        localparam integer d313 = 5;
        for (n313 = 0; n313 < 16; n313 = n313 + 1) 
        begin: outbit313
            assign data_11[n313 + d313*16 + c11*28*16] = data_11_array[c11][d313][n313];
        end
    endgenerate
    generate 
        localparam integer d314 = 6;
        for (n314 = 0; n314 < 16; n314 = n314 + 1) 
        begin: outbit314
            assign data_11[n314 + d314*16 + c11*28*16] = data_11_array[c11][d314][n314];
        end
    endgenerate
    generate 
        localparam integer d315 = 7;
        for (n315 = 0; n315 < 16; n315 = n315 + 1) 
        begin: outbit315
            assign data_11[n315 + d315*16 + c11*28*16] = data_11_array[c11][d315][n315];
        end
    endgenerate
    generate 
        localparam integer d316 = 8;
        for (n316 = 0; n316 < 16; n316 = n316 + 1) 
        begin: outbit316
            assign data_11[n316 + d316*16 + c11*28*16] = data_11_array[c11][d316][n316];
        end
    endgenerate
    generate 
        localparam integer d317 = 9;
        for (n317 = 0; n317 < 16; n317 = n317 + 1) 
        begin: outbit317
            assign data_11[n317 + d317*16 + c11*28*16] = data_11_array[c11][d317][n317];
        end
    endgenerate
    generate 
        localparam integer d318 = 10;
        for (n318 = 0; n318 < 16; n318 = n318 + 1) 
        begin: outbit318
            assign data_11[n318 + d318*16 + c11*28*16] = data_11_array[c11][d318][n318];
        end
    endgenerate
    generate 
        localparam integer d319 = 11;
        for (n319 = 0; n319 < 16; n319 = n319 + 1) 
        begin: outbit319
            assign data_11[n319 + d319*16 + c11*28*16] = data_11_array[c11][d319][n319];
        end
    endgenerate
    generate 
        localparam integer d320 = 12;
        for (n320 = 0; n320 < 16; n320 = n320 + 1) 
        begin: outbit320
            assign data_11[n320 + d320*16 + c11*28*16] = data_11_array[c11][d320][n320];
        end
    endgenerate
    generate 
        localparam integer d321 = 13;
        for (n321 = 0; n321 < 16; n321 = n321 + 1) 
        begin: outbit321
            assign data_11[n321 + d321*16 + c11*28*16] = data_11_array[c11][d321][n321];
        end
    endgenerate
    generate 
        localparam integer d322 = 14;
        for (n322 = 0; n322 < 16; n322 = n322 + 1) 
        begin: outbit322
            assign data_11[n322 + d322*16 + c11*28*16] = data_11_array[c11][d322][n322];
        end
    endgenerate
    generate 
        localparam integer d323 = 15;
        for (n323 = 0; n323 < 16; n323 = n323 + 1) 
        begin: outbit323
            assign data_11[n323 + d323*16 + c11*28*16] = data_11_array[c11][d323][n323];
        end
    endgenerate
    generate 
        localparam integer d324 = 16;
        for (n324 = 0; n324 < 16; n324 = n324 + 1) 
        begin: outbit324
            assign data_11[n324 + d324*16 + c11*28*16] = data_11_array[c11][d324][n324];
        end
    endgenerate
    generate 
        localparam integer d325 = 17;
        for (n325 = 0; n325 < 16; n325 = n325 + 1) 
        begin: outbit325
            assign data_11[n325 + d325*16 + c11*28*16] = data_11_array[c11][d325][n325];
        end
    endgenerate
    generate 
        localparam integer d326 = 18;
        for (n326 = 0; n326 < 16; n326 = n326 + 1) 
        begin: outbit326
            assign data_11[n326 + d326*16 + c11*28*16] = data_11_array[c11][d326][n326];
        end
    endgenerate
    generate 
        localparam integer d327 = 19;
        for (n327 = 0; n327 < 16; n327 = n327 + 1) 
        begin: outbit327
            assign data_11[n327 + d327*16 + c11*28*16] = data_11_array[c11][d327][n327];
        end
    endgenerate
    generate 
        localparam integer d328 = 20;
        for (n328 = 0; n328 < 16; n328 = n328 + 1) 
        begin: outbit328
            assign data_11[n328 + d328*16 + c11*28*16] = data_11_array[c11][d328][n328];
        end
    endgenerate
    generate 
        localparam integer d329 = 21;
        for (n329 = 0; n329 < 16; n329 = n329 + 1) 
        begin: outbit329
            assign data_11[n329 + d329*16 + c11*28*16] = data_11_array[c11][d329][n329];
        end
    endgenerate
    generate 
        localparam integer d330 = 22;
        for (n330 = 0; n330 < 16; n330 = n330 + 1) 
        begin: outbit330
            assign data_11[n330 + d330*16 + c11*28*16] = data_11_array[c11][d330][n330];
        end
    endgenerate
    generate 
        localparam integer d331 = 23;
        for (n331 = 0; n331 < 16; n331 = n331 + 1) 
        begin: outbit331
            assign data_11[n331 + d331*16 + c11*28*16] = data_11_array[c11][d331][n331];
        end
    endgenerate
    generate 
        localparam integer d332 = 24;
        for (n332 = 0; n332 < 16; n332 = n332 + 1) 
        begin: outbit332
            assign data_11[n332 + d332*16 + c11*28*16] = data_11_array[c11][d332][n332];
        end
    endgenerate
    generate 
        localparam integer d333 = 25;
        for (n333 = 0; n333 < 16; n333 = n333 + 1) 
        begin: outbit333
            assign data_11[n333 + d333*16 + c11*28*16] = data_11_array[c11][d333][n333];
        end
    endgenerate
    generate 
        localparam integer d334 = 26;
        for (n334 = 0; n334 < 16; n334 = n334 + 1) 
        begin: outbit334
            assign data_11[n334 + d334*16 + c11*28*16] = data_11_array[c11][d334][n334];
        end
    endgenerate
    generate 
        localparam integer d335 = 27;
        for (n335 = 0; n335 < 16; n335 = n335 + 1) 
        begin: outbit335
            assign data_11[n335 + d335*16 + c11*28*16] = data_11_array[c11][d335][n335];
        end
    endgenerate
    localparam integer c12 = 12;
    generate 
        localparam integer d336 = 0;
        for (n336 = 0; n336 < 16; n336 = n336 + 1) 
        begin: outbit336
            assign data_11[n336 + d336*16 + c12*28*16] = data_11_array[c12][d336][n336];
        end
    endgenerate
    generate 
        localparam integer d337 = 1;
        for (n337 = 0; n337 < 16; n337 = n337 + 1) 
        begin: outbit337
            assign data_11[n337 + d337*16 + c12*28*16] = data_11_array[c12][d337][n337];
        end
    endgenerate
    generate 
        localparam integer d338 = 2;
        for (n338 = 0; n338 < 16; n338 = n338 + 1) 
        begin: outbit338
            assign data_11[n338 + d338*16 + c12*28*16] = data_11_array[c12][d338][n338];
        end
    endgenerate
    generate 
        localparam integer d339 = 3;
        for (n339 = 0; n339 < 16; n339 = n339 + 1) 
        begin: outbit339
            assign data_11[n339 + d339*16 + c12*28*16] = data_11_array[c12][d339][n339];
        end
    endgenerate
    generate 
        localparam integer d340 = 4;
        for (n340 = 0; n340 < 16; n340 = n340 + 1) 
        begin: outbit340
            assign data_11[n340 + d340*16 + c12*28*16] = data_11_array[c12][d340][n340];
        end
    endgenerate
    generate 
        localparam integer d341 = 5;
        for (n341 = 0; n341 < 16; n341 = n341 + 1) 
        begin: outbit341
            assign data_11[n341 + d341*16 + c12*28*16] = data_11_array[c12][d341][n341];
        end
    endgenerate
    generate 
        localparam integer d342 = 6;
        for (n342 = 0; n342 < 16; n342 = n342 + 1) 
        begin: outbit342
            assign data_11[n342 + d342*16 + c12*28*16] = data_11_array[c12][d342][n342];
        end
    endgenerate
    generate 
        localparam integer d343 = 7;
        for (n343 = 0; n343 < 16; n343 = n343 + 1) 
        begin: outbit343
            assign data_11[n343 + d343*16 + c12*28*16] = data_11_array[c12][d343][n343];
        end
    endgenerate
    generate 
        localparam integer d344 = 8;
        for (n344 = 0; n344 < 16; n344 = n344 + 1) 
        begin: outbit344
            assign data_11[n344 + d344*16 + c12*28*16] = data_11_array[c12][d344][n344];
        end
    endgenerate
    generate 
        localparam integer d345 = 9;
        for (n345 = 0; n345 < 16; n345 = n345 + 1) 
        begin: outbit345
            assign data_11[n345 + d345*16 + c12*28*16] = data_11_array[c12][d345][n345];
        end
    endgenerate
    generate 
        localparam integer d346 = 10;
        for (n346 = 0; n346 < 16; n346 = n346 + 1) 
        begin: outbit346
            assign data_11[n346 + d346*16 + c12*28*16] = data_11_array[c12][d346][n346];
        end
    endgenerate
    generate 
        localparam integer d347 = 11;
        for (n347 = 0; n347 < 16; n347 = n347 + 1) 
        begin: outbit347
            assign data_11[n347 + d347*16 + c12*28*16] = data_11_array[c12][d347][n347];
        end
    endgenerate
    generate 
        localparam integer d348 = 12;
        for (n348 = 0; n348 < 16; n348 = n348 + 1) 
        begin: outbit348
            assign data_11[n348 + d348*16 + c12*28*16] = data_11_array[c12][d348][n348];
        end
    endgenerate
    generate 
        localparam integer d349 = 13;
        for (n349 = 0; n349 < 16; n349 = n349 + 1) 
        begin: outbit349
            assign data_11[n349 + d349*16 + c12*28*16] = data_11_array[c12][d349][n349];
        end
    endgenerate
    generate 
        localparam integer d350 = 14;
        for (n350 = 0; n350 < 16; n350 = n350 + 1) 
        begin: outbit350
            assign data_11[n350 + d350*16 + c12*28*16] = data_11_array[c12][d350][n350];
        end
    endgenerate
    generate 
        localparam integer d351 = 15;
        for (n351 = 0; n351 < 16; n351 = n351 + 1) 
        begin: outbit351
            assign data_11[n351 + d351*16 + c12*28*16] = data_11_array[c12][d351][n351];
        end
    endgenerate
    generate 
        localparam integer d352 = 16;
        for (n352 = 0; n352 < 16; n352 = n352 + 1) 
        begin: outbit352
            assign data_11[n352 + d352*16 + c12*28*16] = data_11_array[c12][d352][n352];
        end
    endgenerate
    generate 
        localparam integer d353 = 17;
        for (n353 = 0; n353 < 16; n353 = n353 + 1) 
        begin: outbit353
            assign data_11[n353 + d353*16 + c12*28*16] = data_11_array[c12][d353][n353];
        end
    endgenerate
    generate 
        localparam integer d354 = 18;
        for (n354 = 0; n354 < 16; n354 = n354 + 1) 
        begin: outbit354
            assign data_11[n354 + d354*16 + c12*28*16] = data_11_array[c12][d354][n354];
        end
    endgenerate
    generate 
        localparam integer d355 = 19;
        for (n355 = 0; n355 < 16; n355 = n355 + 1) 
        begin: outbit355
            assign data_11[n355 + d355*16 + c12*28*16] = data_11_array[c12][d355][n355];
        end
    endgenerate
    generate 
        localparam integer d356 = 20;
        for (n356 = 0; n356 < 16; n356 = n356 + 1) 
        begin: outbit356
            assign data_11[n356 + d356*16 + c12*28*16] = data_11_array[c12][d356][n356];
        end
    endgenerate
    generate 
        localparam integer d357 = 21;
        for (n357 = 0; n357 < 16; n357 = n357 + 1) 
        begin: outbit357
            assign data_11[n357 + d357*16 + c12*28*16] = data_11_array[c12][d357][n357];
        end
    endgenerate
    generate 
        localparam integer d358 = 22;
        for (n358 = 0; n358 < 16; n358 = n358 + 1) 
        begin: outbit358
            assign data_11[n358 + d358*16 + c12*28*16] = data_11_array[c12][d358][n358];
        end
    endgenerate
    generate 
        localparam integer d359 = 23;
        for (n359 = 0; n359 < 16; n359 = n359 + 1) 
        begin: outbit359
            assign data_11[n359 + d359*16 + c12*28*16] = data_11_array[c12][d359][n359];
        end
    endgenerate
    generate 
        localparam integer d360 = 24;
        for (n360 = 0; n360 < 16; n360 = n360 + 1) 
        begin: outbit360
            assign data_11[n360 + d360*16 + c12*28*16] = data_11_array[c12][d360][n360];
        end
    endgenerate
    generate 
        localparam integer d361 = 25;
        for (n361 = 0; n361 < 16; n361 = n361 + 1) 
        begin: outbit361
            assign data_11[n361 + d361*16 + c12*28*16] = data_11_array[c12][d361][n361];
        end
    endgenerate
    generate 
        localparam integer d362 = 26;
        for (n362 = 0; n362 < 16; n362 = n362 + 1) 
        begin: outbit362
            assign data_11[n362 + d362*16 + c12*28*16] = data_11_array[c12][d362][n362];
        end
    endgenerate
    generate 
        localparam integer d363 = 27;
        for (n363 = 0; n363 < 16; n363 = n363 + 1) 
        begin: outbit363
            assign data_11[n363 + d363*16 + c12*28*16] = data_11_array[c12][d363][n363];
        end
    endgenerate
    localparam integer c13 = 13;
    generate 
        localparam integer d364 = 0;
        for (n364 = 0; n364 < 16; n364 = n364 + 1) 
        begin: outbit364
            assign data_11[n364 + d364*16 + c13*28*16] = data_11_array[c13][d364][n364];
        end
    endgenerate
    generate 
        localparam integer d365 = 1;
        for (n365 = 0; n365 < 16; n365 = n365 + 1) 
        begin: outbit365
            assign data_11[n365 + d365*16 + c13*28*16] = data_11_array[c13][d365][n365];
        end
    endgenerate
    generate 
        localparam integer d366 = 2;
        for (n366 = 0; n366 < 16; n366 = n366 + 1) 
        begin: outbit366
            assign data_11[n366 + d366*16 + c13*28*16] = data_11_array[c13][d366][n366];
        end
    endgenerate
    generate 
        localparam integer d367 = 3;
        for (n367 = 0; n367 < 16; n367 = n367 + 1) 
        begin: outbit367
            assign data_11[n367 + d367*16 + c13*28*16] = data_11_array[c13][d367][n367];
        end
    endgenerate
    generate 
        localparam integer d368 = 4;
        for (n368 = 0; n368 < 16; n368 = n368 + 1) 
        begin: outbit368
            assign data_11[n368 + d368*16 + c13*28*16] = data_11_array[c13][d368][n368];
        end
    endgenerate
    generate 
        localparam integer d369 = 5;
        for (n369 = 0; n369 < 16; n369 = n369 + 1) 
        begin: outbit369
            assign data_11[n369 + d369*16 + c13*28*16] = data_11_array[c13][d369][n369];
        end
    endgenerate
    generate 
        localparam integer d370 = 6;
        for (n370 = 0; n370 < 16; n370 = n370 + 1) 
        begin: outbit370
            assign data_11[n370 + d370*16 + c13*28*16] = data_11_array[c13][d370][n370];
        end
    endgenerate
    generate 
        localparam integer d371 = 7;
        for (n371 = 0; n371 < 16; n371 = n371 + 1) 
        begin: outbit371
            assign data_11[n371 + d371*16 + c13*28*16] = data_11_array[c13][d371][n371];
        end
    endgenerate
    generate 
        localparam integer d372 = 8;
        for (n372 = 0; n372 < 16; n372 = n372 + 1) 
        begin: outbit372
            assign data_11[n372 + d372*16 + c13*28*16] = data_11_array[c13][d372][n372];
        end
    endgenerate
    generate 
        localparam integer d373 = 9;
        for (n373 = 0; n373 < 16; n373 = n373 + 1) 
        begin: outbit373
            assign data_11[n373 + d373*16 + c13*28*16] = data_11_array[c13][d373][n373];
        end
    endgenerate
    generate 
        localparam integer d374 = 10;
        for (n374 = 0; n374 < 16; n374 = n374 + 1) 
        begin: outbit374
            assign data_11[n374 + d374*16 + c13*28*16] = data_11_array[c13][d374][n374];
        end
    endgenerate
    generate 
        localparam integer d375 = 11;
        for (n375 = 0; n375 < 16; n375 = n375 + 1) 
        begin: outbit375
            assign data_11[n375 + d375*16 + c13*28*16] = data_11_array[c13][d375][n375];
        end
    endgenerate
    generate 
        localparam integer d376 = 12;
        for (n376 = 0; n376 < 16; n376 = n376 + 1) 
        begin: outbit376
            assign data_11[n376 + d376*16 + c13*28*16] = data_11_array[c13][d376][n376];
        end
    endgenerate
    generate 
        localparam integer d377 = 13;
        for (n377 = 0; n377 < 16; n377 = n377 + 1) 
        begin: outbit377
            assign data_11[n377 + d377*16 + c13*28*16] = data_11_array[c13][d377][n377];
        end
    endgenerate
    generate 
        localparam integer d378 = 14;
        for (n378 = 0; n378 < 16; n378 = n378 + 1) 
        begin: outbit378
            assign data_11[n378 + d378*16 + c13*28*16] = data_11_array[c13][d378][n378];
        end
    endgenerate
    generate 
        localparam integer d379 = 15;
        for (n379 = 0; n379 < 16; n379 = n379 + 1) 
        begin: outbit379
            assign data_11[n379 + d379*16 + c13*28*16] = data_11_array[c13][d379][n379];
        end
    endgenerate
    generate 
        localparam integer d380 = 16;
        for (n380 = 0; n380 < 16; n380 = n380 + 1) 
        begin: outbit380
            assign data_11[n380 + d380*16 + c13*28*16] = data_11_array[c13][d380][n380];
        end
    endgenerate
    generate 
        localparam integer d381 = 17;
        for (n381 = 0; n381 < 16; n381 = n381 + 1) 
        begin: outbit381
            assign data_11[n381 + d381*16 + c13*28*16] = data_11_array[c13][d381][n381];
        end
    endgenerate
    generate 
        localparam integer d382 = 18;
        for (n382 = 0; n382 < 16; n382 = n382 + 1) 
        begin: outbit382
            assign data_11[n382 + d382*16 + c13*28*16] = data_11_array[c13][d382][n382];
        end
    endgenerate
    generate 
        localparam integer d383 = 19;
        for (n383 = 0; n383 < 16; n383 = n383 + 1) 
        begin: outbit383
            assign data_11[n383 + d383*16 + c13*28*16] = data_11_array[c13][d383][n383];
        end
    endgenerate
    generate 
        localparam integer d384 = 20;
        for (n384 = 0; n384 < 16; n384 = n384 + 1) 
        begin: outbit384
            assign data_11[n384 + d384*16 + c13*28*16] = data_11_array[c13][d384][n384];
        end
    endgenerate
    generate 
        localparam integer d385 = 21;
        for (n385 = 0; n385 < 16; n385 = n385 + 1) 
        begin: outbit385
            assign data_11[n385 + d385*16 + c13*28*16] = data_11_array[c13][d385][n385];
        end
    endgenerate
    generate 
        localparam integer d386 = 22;
        for (n386 = 0; n386 < 16; n386 = n386 + 1) 
        begin: outbit386
            assign data_11[n386 + d386*16 + c13*28*16] = data_11_array[c13][d386][n386];
        end
    endgenerate
    generate 
        localparam integer d387 = 23;
        for (n387 = 0; n387 < 16; n387 = n387 + 1) 
        begin: outbit387
            assign data_11[n387 + d387*16 + c13*28*16] = data_11_array[c13][d387][n387];
        end
    endgenerate
    generate 
        localparam integer d388 = 24;
        for (n388 = 0; n388 < 16; n388 = n388 + 1) 
        begin: outbit388
            assign data_11[n388 + d388*16 + c13*28*16] = data_11_array[c13][d388][n388];
        end
    endgenerate
    generate 
        localparam integer d389 = 25;
        for (n389 = 0; n389 < 16; n389 = n389 + 1) 
        begin: outbit389
            assign data_11[n389 + d389*16 + c13*28*16] = data_11_array[c13][d389][n389];
        end
    endgenerate
    generate 
        localparam integer d390 = 26;
        for (n390 = 0; n390 < 16; n390 = n390 + 1) 
        begin: outbit390
            assign data_11[n390 + d390*16 + c13*28*16] = data_11_array[c13][d390][n390];
        end
    endgenerate
    generate 
        localparam integer d391 = 27;
        for (n391 = 0; n391 < 16; n391 = n391 + 1) 
        begin: outbit391
            assign data_11[n391 + d391*16 + c13*28*16] = data_11_array[c13][d391][n391];
        end
    endgenerate
    localparam integer c14 = 14;
    generate 
        localparam integer d392 = 0;
        for (n392 = 0; n392 < 16; n392 = n392 + 1) 
        begin: outbit392
            assign data_11[n392 + d392*16 + c14*28*16] = data_11_array[c14][d392][n392];
        end
    endgenerate
    generate 
        localparam integer d393 = 1;
        for (n393 = 0; n393 < 16; n393 = n393 + 1) 
        begin: outbit393
            assign data_11[n393 + d393*16 + c14*28*16] = data_11_array[c14][d393][n393];
        end
    endgenerate
    generate 
        localparam integer d394 = 2;
        for (n394 = 0; n394 < 16; n394 = n394 + 1) 
        begin: outbit394
            assign data_11[n394 + d394*16 + c14*28*16] = data_11_array[c14][d394][n394];
        end
    endgenerate
    generate 
        localparam integer d395 = 3;
        for (n395 = 0; n395 < 16; n395 = n395 + 1) 
        begin: outbit395
            assign data_11[n395 + d395*16 + c14*28*16] = data_11_array[c14][d395][n395];
        end
    endgenerate
    generate 
        localparam integer d396 = 4;
        for (n396 = 0; n396 < 16; n396 = n396 + 1) 
        begin: outbit396
            assign data_11[n396 + d396*16 + c14*28*16] = data_11_array[c14][d396][n396];
        end
    endgenerate
    generate 
        localparam integer d397 = 5;
        for (n397 = 0; n397 < 16; n397 = n397 + 1) 
        begin: outbit397
            assign data_11[n397 + d397*16 + c14*28*16] = data_11_array[c14][d397][n397];
        end
    endgenerate
    generate 
        localparam integer d398 = 6;
        for (n398 = 0; n398 < 16; n398 = n398 + 1) 
        begin: outbit398
            assign data_11[n398 + d398*16 + c14*28*16] = data_11_array[c14][d398][n398];
        end
    endgenerate
    generate 
        localparam integer d399 = 7;
        for (n399 = 0; n399 < 16; n399 = n399 + 1) 
        begin: outbit399
            assign data_11[n399 + d399*16 + c14*28*16] = data_11_array[c14][d399][n399];
        end
    endgenerate
    generate 
        localparam integer d400 = 8;
        for (n400 = 0; n400 < 16; n400 = n400 + 1) 
        begin: outbit400
            assign data_11[n400 + d400*16 + c14*28*16] = data_11_array[c14][d400][n400];
        end
    endgenerate
    generate 
        localparam integer d401 = 9;
        for (n401 = 0; n401 < 16; n401 = n401 + 1) 
        begin: outbit401
            assign data_11[n401 + d401*16 + c14*28*16] = data_11_array[c14][d401][n401];
        end
    endgenerate
    generate 
        localparam integer d402 = 10;
        for (n402 = 0; n402 < 16; n402 = n402 + 1) 
        begin: outbit402
            assign data_11[n402 + d402*16 + c14*28*16] = data_11_array[c14][d402][n402];
        end
    endgenerate
    generate 
        localparam integer d403 = 11;
        for (n403 = 0; n403 < 16; n403 = n403 + 1) 
        begin: outbit403
            assign data_11[n403 + d403*16 + c14*28*16] = data_11_array[c14][d403][n403];
        end
    endgenerate
    generate 
        localparam integer d404 = 12;
        for (n404 = 0; n404 < 16; n404 = n404 + 1) 
        begin: outbit404
            assign data_11[n404 + d404*16 + c14*28*16] = data_11_array[c14][d404][n404];
        end
    endgenerate
    generate 
        localparam integer d405 = 13;
        for (n405 = 0; n405 < 16; n405 = n405 + 1) 
        begin: outbit405
            assign data_11[n405 + d405*16 + c14*28*16] = data_11_array[c14][d405][n405];
        end
    endgenerate
    generate 
        localparam integer d406 = 14;
        for (n406 = 0; n406 < 16; n406 = n406 + 1) 
        begin: outbit406
            assign data_11[n406 + d406*16 + c14*28*16] = data_11_array[c14][d406][n406];
        end
    endgenerate
    generate 
        localparam integer d407 = 15;
        for (n407 = 0; n407 < 16; n407 = n407 + 1) 
        begin: outbit407
            assign data_11[n407 + d407*16 + c14*28*16] = data_11_array[c14][d407][n407];
        end
    endgenerate
    generate 
        localparam integer d408 = 16;
        for (n408 = 0; n408 < 16; n408 = n408 + 1) 
        begin: outbit408
            assign data_11[n408 + d408*16 + c14*28*16] = data_11_array[c14][d408][n408];
        end
    endgenerate
    generate 
        localparam integer d409 = 17;
        for (n409 = 0; n409 < 16; n409 = n409 + 1) 
        begin: outbit409
            assign data_11[n409 + d409*16 + c14*28*16] = data_11_array[c14][d409][n409];
        end
    endgenerate
    generate 
        localparam integer d410 = 18;
        for (n410 = 0; n410 < 16; n410 = n410 + 1) 
        begin: outbit410
            assign data_11[n410 + d410*16 + c14*28*16] = data_11_array[c14][d410][n410];
        end
    endgenerate
    generate 
        localparam integer d411 = 19;
        for (n411 = 0; n411 < 16; n411 = n411 + 1) 
        begin: outbit411
            assign data_11[n411 + d411*16 + c14*28*16] = data_11_array[c14][d411][n411];
        end
    endgenerate
    generate 
        localparam integer d412 = 20;
        for (n412 = 0; n412 < 16; n412 = n412 + 1) 
        begin: outbit412
            assign data_11[n412 + d412*16 + c14*28*16] = data_11_array[c14][d412][n412];
        end
    endgenerate
    generate 
        localparam integer d413 = 21;
        for (n413 = 0; n413 < 16; n413 = n413 + 1) 
        begin: outbit413
            assign data_11[n413 + d413*16 + c14*28*16] = data_11_array[c14][d413][n413];
        end
    endgenerate
    generate 
        localparam integer d414 = 22;
        for (n414 = 0; n414 < 16; n414 = n414 + 1) 
        begin: outbit414
            assign data_11[n414 + d414*16 + c14*28*16] = data_11_array[c14][d414][n414];
        end
    endgenerate
    generate 
        localparam integer d415 = 23;
        for (n415 = 0; n415 < 16; n415 = n415 + 1) 
        begin: outbit415
            assign data_11[n415 + d415*16 + c14*28*16] = data_11_array[c14][d415][n415];
        end
    endgenerate
    generate 
        localparam integer d416 = 24;
        for (n416 = 0; n416 < 16; n416 = n416 + 1) 
        begin: outbit416
            assign data_11[n416 + d416*16 + c14*28*16] = data_11_array[c14][d416][n416];
        end
    endgenerate
    generate 
        localparam integer d417 = 25;
        for (n417 = 0; n417 < 16; n417 = n417 + 1) 
        begin: outbit417
            assign data_11[n417 + d417*16 + c14*28*16] = data_11_array[c14][d417][n417];
        end
    endgenerate
    generate 
        localparam integer d418 = 26;
        for (n418 = 0; n418 < 16; n418 = n418 + 1) 
        begin: outbit418
            assign data_11[n418 + d418*16 + c14*28*16] = data_11_array[c14][d418][n418];
        end
    endgenerate
    generate 
        localparam integer d419 = 27;
        for (n419 = 0; n419 < 16; n419 = n419 + 1) 
        begin: outbit419
            assign data_11[n419 + d419*16 + c14*28*16] = data_11_array[c14][d419][n419];
        end
    endgenerate
    localparam integer c15 = 15;
    generate 
        localparam integer d420 = 0;
        for (n420 = 0; n420 < 16; n420 = n420 + 1) 
        begin: outbit420
            assign data_11[n420 + d420*16 + c15*28*16] = data_11_array[c15][d420][n420];
        end
    endgenerate
    generate 
        localparam integer d421 = 1;
        for (n421 = 0; n421 < 16; n421 = n421 + 1) 
        begin: outbit421
            assign data_11[n421 + d421*16 + c15*28*16] = data_11_array[c15][d421][n421];
        end
    endgenerate
    generate 
        localparam integer d422 = 2;
        for (n422 = 0; n422 < 16; n422 = n422 + 1) 
        begin: outbit422
            assign data_11[n422 + d422*16 + c15*28*16] = data_11_array[c15][d422][n422];
        end
    endgenerate
    generate 
        localparam integer d423 = 3;
        for (n423 = 0; n423 < 16; n423 = n423 + 1) 
        begin: outbit423
            assign data_11[n423 + d423*16 + c15*28*16] = data_11_array[c15][d423][n423];
        end
    endgenerate
    generate 
        localparam integer d424 = 4;
        for (n424 = 0; n424 < 16; n424 = n424 + 1) 
        begin: outbit424
            assign data_11[n424 + d424*16 + c15*28*16] = data_11_array[c15][d424][n424];
        end
    endgenerate
    generate 
        localparam integer d425 = 5;
        for (n425 = 0; n425 < 16; n425 = n425 + 1) 
        begin: outbit425
            assign data_11[n425 + d425*16 + c15*28*16] = data_11_array[c15][d425][n425];
        end
    endgenerate
    generate 
        localparam integer d426 = 6;
        for (n426 = 0; n426 < 16; n426 = n426 + 1) 
        begin: outbit426
            assign data_11[n426 + d426*16 + c15*28*16] = data_11_array[c15][d426][n426];
        end
    endgenerate
    generate 
        localparam integer d427 = 7;
        for (n427 = 0; n427 < 16; n427 = n427 + 1) 
        begin: outbit427
            assign data_11[n427 + d427*16 + c15*28*16] = data_11_array[c15][d427][n427];
        end
    endgenerate
    generate 
        localparam integer d428 = 8;
        for (n428 = 0; n428 < 16; n428 = n428 + 1) 
        begin: outbit428
            assign data_11[n428 + d428*16 + c15*28*16] = data_11_array[c15][d428][n428];
        end
    endgenerate
    generate 
        localparam integer d429 = 9;
        for (n429 = 0; n429 < 16; n429 = n429 + 1) 
        begin: outbit429
            assign data_11[n429 + d429*16 + c15*28*16] = data_11_array[c15][d429][n429];
        end
    endgenerate
    generate 
        localparam integer d430 = 10;
        for (n430 = 0; n430 < 16; n430 = n430 + 1) 
        begin: outbit430
            assign data_11[n430 + d430*16 + c15*28*16] = data_11_array[c15][d430][n430];
        end
    endgenerate
    generate 
        localparam integer d431 = 11;
        for (n431 = 0; n431 < 16; n431 = n431 + 1) 
        begin: outbit431
            assign data_11[n431 + d431*16 + c15*28*16] = data_11_array[c15][d431][n431];
        end
    endgenerate
    generate 
        localparam integer d432 = 12;
        for (n432 = 0; n432 < 16; n432 = n432 + 1) 
        begin: outbit432
            assign data_11[n432 + d432*16 + c15*28*16] = data_11_array[c15][d432][n432];
        end
    endgenerate
    generate 
        localparam integer d433 = 13;
        for (n433 = 0; n433 < 16; n433 = n433 + 1) 
        begin: outbit433
            assign data_11[n433 + d433*16 + c15*28*16] = data_11_array[c15][d433][n433];
        end
    endgenerate
    generate 
        localparam integer d434 = 14;
        for (n434 = 0; n434 < 16; n434 = n434 + 1) 
        begin: outbit434
            assign data_11[n434 + d434*16 + c15*28*16] = data_11_array[c15][d434][n434];
        end
    endgenerate
    generate 
        localparam integer d435 = 15;
        for (n435 = 0; n435 < 16; n435 = n435 + 1) 
        begin: outbit435
            assign data_11[n435 + d435*16 + c15*28*16] = data_11_array[c15][d435][n435];
        end
    endgenerate
    generate 
        localparam integer d436 = 16;
        for (n436 = 0; n436 < 16; n436 = n436 + 1) 
        begin: outbit436
            assign data_11[n436 + d436*16 + c15*28*16] = data_11_array[c15][d436][n436];
        end
    endgenerate
    generate 
        localparam integer d437 = 17;
        for (n437 = 0; n437 < 16; n437 = n437 + 1) 
        begin: outbit437
            assign data_11[n437 + d437*16 + c15*28*16] = data_11_array[c15][d437][n437];
        end
    endgenerate
    generate 
        localparam integer d438 = 18;
        for (n438 = 0; n438 < 16; n438 = n438 + 1) 
        begin: outbit438
            assign data_11[n438 + d438*16 + c15*28*16] = data_11_array[c15][d438][n438];
        end
    endgenerate
    generate 
        localparam integer d439 = 19;
        for (n439 = 0; n439 < 16; n439 = n439 + 1) 
        begin: outbit439
            assign data_11[n439 + d439*16 + c15*28*16] = data_11_array[c15][d439][n439];
        end
    endgenerate
    generate 
        localparam integer d440 = 20;
        for (n440 = 0; n440 < 16; n440 = n440 + 1) 
        begin: outbit440
            assign data_11[n440 + d440*16 + c15*28*16] = data_11_array[c15][d440][n440];
        end
    endgenerate
    generate 
        localparam integer d441 = 21;
        for (n441 = 0; n441 < 16; n441 = n441 + 1) 
        begin: outbit441
            assign data_11[n441 + d441*16 + c15*28*16] = data_11_array[c15][d441][n441];
        end
    endgenerate
    generate 
        localparam integer d442 = 22;
        for (n442 = 0; n442 < 16; n442 = n442 + 1) 
        begin: outbit442
            assign data_11[n442 + d442*16 + c15*28*16] = data_11_array[c15][d442][n442];
        end
    endgenerate
    generate 
        localparam integer d443 = 23;
        for (n443 = 0; n443 < 16; n443 = n443 + 1) 
        begin: outbit443
            assign data_11[n443 + d443*16 + c15*28*16] = data_11_array[c15][d443][n443];
        end
    endgenerate
    generate 
        localparam integer d444 = 24;
        for (n444 = 0; n444 < 16; n444 = n444 + 1) 
        begin: outbit444
            assign data_11[n444 + d444*16 + c15*28*16] = data_11_array[c15][d444][n444];
        end
    endgenerate
    generate 
        localparam integer d445 = 25;
        for (n445 = 0; n445 < 16; n445 = n445 + 1) 
        begin: outbit445
            assign data_11[n445 + d445*16 + c15*28*16] = data_11_array[c15][d445][n445];
        end
    endgenerate
    generate 
        localparam integer d446 = 26;
        for (n446 = 0; n446 < 16; n446 = n446 + 1) 
        begin: outbit446
            assign data_11[n446 + d446*16 + c15*28*16] = data_11_array[c15][d446][n446];
        end
    endgenerate
    generate 
        localparam integer d447 = 27;
        for (n447 = 0; n447 < 16; n447 = n447 + 1) 
        begin: outbit447
            assign data_11[n447 + d447*16 + c15*28*16] = data_11_array[c15][d447][n447];
        end
    endgenerate
    localparam integer c16 = 16;
    generate 
        localparam integer d448 = 0;
        for (n448 = 0; n448 < 16; n448 = n448 + 1) 
        begin: outbit448
            assign data_11[n448 + d448*16 + c16*28*16] = data_11_array[c16][d448][n448];
        end
    endgenerate
    generate 
        localparam integer d449 = 1;
        for (n449 = 0; n449 < 16; n449 = n449 + 1) 
        begin: outbit449
            assign data_11[n449 + d449*16 + c16*28*16] = data_11_array[c16][d449][n449];
        end
    endgenerate
    generate 
        localparam integer d450 = 2;
        for (n450 = 0; n450 < 16; n450 = n450 + 1) 
        begin: outbit450
            assign data_11[n450 + d450*16 + c16*28*16] = data_11_array[c16][d450][n450];
        end
    endgenerate
    generate 
        localparam integer d451 = 3;
        for (n451 = 0; n451 < 16; n451 = n451 + 1) 
        begin: outbit451
            assign data_11[n451 + d451*16 + c16*28*16] = data_11_array[c16][d451][n451];
        end
    endgenerate
    generate 
        localparam integer d452 = 4;
        for (n452 = 0; n452 < 16; n452 = n452 + 1) 
        begin: outbit452
            assign data_11[n452 + d452*16 + c16*28*16] = data_11_array[c16][d452][n452];
        end
    endgenerate
    generate 
        localparam integer d453 = 5;
        for (n453 = 0; n453 < 16; n453 = n453 + 1) 
        begin: outbit453
            assign data_11[n453 + d453*16 + c16*28*16] = data_11_array[c16][d453][n453];
        end
    endgenerate
    generate 
        localparam integer d454 = 6;
        for (n454 = 0; n454 < 16; n454 = n454 + 1) 
        begin: outbit454
            assign data_11[n454 + d454*16 + c16*28*16] = data_11_array[c16][d454][n454];
        end
    endgenerate
    generate 
        localparam integer d455 = 7;
        for (n455 = 0; n455 < 16; n455 = n455 + 1) 
        begin: outbit455
            assign data_11[n455 + d455*16 + c16*28*16] = data_11_array[c16][d455][n455];
        end
    endgenerate
    generate 
        localparam integer d456 = 8;
        for (n456 = 0; n456 < 16; n456 = n456 + 1) 
        begin: outbit456
            assign data_11[n456 + d456*16 + c16*28*16] = data_11_array[c16][d456][n456];
        end
    endgenerate
    generate 
        localparam integer d457 = 9;
        for (n457 = 0; n457 < 16; n457 = n457 + 1) 
        begin: outbit457
            assign data_11[n457 + d457*16 + c16*28*16] = data_11_array[c16][d457][n457];
        end
    endgenerate
    generate 
        localparam integer d458 = 10;
        for (n458 = 0; n458 < 16; n458 = n458 + 1) 
        begin: outbit458
            assign data_11[n458 + d458*16 + c16*28*16] = data_11_array[c16][d458][n458];
        end
    endgenerate
    generate 
        localparam integer d459 = 11;
        for (n459 = 0; n459 < 16; n459 = n459 + 1) 
        begin: outbit459
            assign data_11[n459 + d459*16 + c16*28*16] = data_11_array[c16][d459][n459];
        end
    endgenerate
    generate 
        localparam integer d460 = 12;
        for (n460 = 0; n460 < 16; n460 = n460 + 1) 
        begin: outbit460
            assign data_11[n460 + d460*16 + c16*28*16] = data_11_array[c16][d460][n460];
        end
    endgenerate
    generate 
        localparam integer d461 = 13;
        for (n461 = 0; n461 < 16; n461 = n461 + 1) 
        begin: outbit461
            assign data_11[n461 + d461*16 + c16*28*16] = data_11_array[c16][d461][n461];
        end
    endgenerate
    generate 
        localparam integer d462 = 14;
        for (n462 = 0; n462 < 16; n462 = n462 + 1) 
        begin: outbit462
            assign data_11[n462 + d462*16 + c16*28*16] = data_11_array[c16][d462][n462];
        end
    endgenerate
    generate 
        localparam integer d463 = 15;
        for (n463 = 0; n463 < 16; n463 = n463 + 1) 
        begin: outbit463
            assign data_11[n463 + d463*16 + c16*28*16] = data_11_array[c16][d463][n463];
        end
    endgenerate
    generate 
        localparam integer d464 = 16;
        for (n464 = 0; n464 < 16; n464 = n464 + 1) 
        begin: outbit464
            assign data_11[n464 + d464*16 + c16*28*16] = data_11_array[c16][d464][n464];
        end
    endgenerate
    generate 
        localparam integer d465 = 17;
        for (n465 = 0; n465 < 16; n465 = n465 + 1) 
        begin: outbit465
            assign data_11[n465 + d465*16 + c16*28*16] = data_11_array[c16][d465][n465];
        end
    endgenerate
    generate 
        localparam integer d466 = 18;
        for (n466 = 0; n466 < 16; n466 = n466 + 1) 
        begin: outbit466
            assign data_11[n466 + d466*16 + c16*28*16] = data_11_array[c16][d466][n466];
        end
    endgenerate
    generate 
        localparam integer d467 = 19;
        for (n467 = 0; n467 < 16; n467 = n467 + 1) 
        begin: outbit467
            assign data_11[n467 + d467*16 + c16*28*16] = data_11_array[c16][d467][n467];
        end
    endgenerate
    generate 
        localparam integer d468 = 20;
        for (n468 = 0; n468 < 16; n468 = n468 + 1) 
        begin: outbit468
            assign data_11[n468 + d468*16 + c16*28*16] = data_11_array[c16][d468][n468];
        end
    endgenerate
    generate 
        localparam integer d469 = 21;
        for (n469 = 0; n469 < 16; n469 = n469 + 1) 
        begin: outbit469
            assign data_11[n469 + d469*16 + c16*28*16] = data_11_array[c16][d469][n469];
        end
    endgenerate
    generate 
        localparam integer d470 = 22;
        for (n470 = 0; n470 < 16; n470 = n470 + 1) 
        begin: outbit470
            assign data_11[n470 + d470*16 + c16*28*16] = data_11_array[c16][d470][n470];
        end
    endgenerate
    generate 
        localparam integer d471 = 23;
        for (n471 = 0; n471 < 16; n471 = n471 + 1) 
        begin: outbit471
            assign data_11[n471 + d471*16 + c16*28*16] = data_11_array[c16][d471][n471];
        end
    endgenerate
    generate 
        localparam integer d472 = 24;
        for (n472 = 0; n472 < 16; n472 = n472 + 1) 
        begin: outbit472
            assign data_11[n472 + d472*16 + c16*28*16] = data_11_array[c16][d472][n472];
        end
    endgenerate
    generate 
        localparam integer d473 = 25;
        for (n473 = 0; n473 < 16; n473 = n473 + 1) 
        begin: outbit473
            assign data_11[n473 + d473*16 + c16*28*16] = data_11_array[c16][d473][n473];
        end
    endgenerate
    generate 
        localparam integer d474 = 26;
        for (n474 = 0; n474 < 16; n474 = n474 + 1) 
        begin: outbit474
            assign data_11[n474 + d474*16 + c16*28*16] = data_11_array[c16][d474][n474];
        end
    endgenerate
    generate 
        localparam integer d475 = 27;
        for (n475 = 0; n475 < 16; n475 = n475 + 1) 
        begin: outbit475
            assign data_11[n475 + d475*16 + c16*28*16] = data_11_array[c16][d475][n475];
        end
    endgenerate
    localparam integer c17 = 17;
    generate 
        localparam integer d476 = 0;
        for (n476 = 0; n476 < 16; n476 = n476 + 1) 
        begin: outbit476
            assign data_11[n476 + d476*16 + c17*28*16] = data_11_array[c17][d476][n476];
        end
    endgenerate
    generate 
        localparam integer d477 = 1;
        for (n477 = 0; n477 < 16; n477 = n477 + 1) 
        begin: outbit477
            assign data_11[n477 + d477*16 + c17*28*16] = data_11_array[c17][d477][n477];
        end
    endgenerate
    generate 
        localparam integer d478 = 2;
        for (n478 = 0; n478 < 16; n478 = n478 + 1) 
        begin: outbit478
            assign data_11[n478 + d478*16 + c17*28*16] = data_11_array[c17][d478][n478];
        end
    endgenerate
    generate 
        localparam integer d479 = 3;
        for (n479 = 0; n479 < 16; n479 = n479 + 1) 
        begin: outbit479
            assign data_11[n479 + d479*16 + c17*28*16] = data_11_array[c17][d479][n479];
        end
    endgenerate
    generate 
        localparam integer d480 = 4;
        for (n480 = 0; n480 < 16; n480 = n480 + 1) 
        begin: outbit480
            assign data_11[n480 + d480*16 + c17*28*16] = data_11_array[c17][d480][n480];
        end
    endgenerate
    generate 
        localparam integer d481 = 5;
        for (n481 = 0; n481 < 16; n481 = n481 + 1) 
        begin: outbit481
            assign data_11[n481 + d481*16 + c17*28*16] = data_11_array[c17][d481][n481];
        end
    endgenerate
    generate 
        localparam integer d482 = 6;
        for (n482 = 0; n482 < 16; n482 = n482 + 1) 
        begin: outbit482
            assign data_11[n482 + d482*16 + c17*28*16] = data_11_array[c17][d482][n482];
        end
    endgenerate
    generate 
        localparam integer d483 = 7;
        for (n483 = 0; n483 < 16; n483 = n483 + 1) 
        begin: outbit483
            assign data_11[n483 + d483*16 + c17*28*16] = data_11_array[c17][d483][n483];
        end
    endgenerate
    generate 
        localparam integer d484 = 8;
        for (n484 = 0; n484 < 16; n484 = n484 + 1) 
        begin: outbit484
            assign data_11[n484 + d484*16 + c17*28*16] = data_11_array[c17][d484][n484];
        end
    endgenerate
    generate 
        localparam integer d485 = 9;
        for (n485 = 0; n485 < 16; n485 = n485 + 1) 
        begin: outbit485
            assign data_11[n485 + d485*16 + c17*28*16] = data_11_array[c17][d485][n485];
        end
    endgenerate
    generate 
        localparam integer d486 = 10;
        for (n486 = 0; n486 < 16; n486 = n486 + 1) 
        begin: outbit486
            assign data_11[n486 + d486*16 + c17*28*16] = data_11_array[c17][d486][n486];
        end
    endgenerate
    generate 
        localparam integer d487 = 11;
        for (n487 = 0; n487 < 16; n487 = n487 + 1) 
        begin: outbit487
            assign data_11[n487 + d487*16 + c17*28*16] = data_11_array[c17][d487][n487];
        end
    endgenerate
    generate 
        localparam integer d488 = 12;
        for (n488 = 0; n488 < 16; n488 = n488 + 1) 
        begin: outbit488
            assign data_11[n488 + d488*16 + c17*28*16] = data_11_array[c17][d488][n488];
        end
    endgenerate
    generate 
        localparam integer d489 = 13;
        for (n489 = 0; n489 < 16; n489 = n489 + 1) 
        begin: outbit489
            assign data_11[n489 + d489*16 + c17*28*16] = data_11_array[c17][d489][n489];
        end
    endgenerate
    generate 
        localparam integer d490 = 14;
        for (n490 = 0; n490 < 16; n490 = n490 + 1) 
        begin: outbit490
            assign data_11[n490 + d490*16 + c17*28*16] = data_11_array[c17][d490][n490];
        end
    endgenerate
    generate 
        localparam integer d491 = 15;
        for (n491 = 0; n491 < 16; n491 = n491 + 1) 
        begin: outbit491
            assign data_11[n491 + d491*16 + c17*28*16] = data_11_array[c17][d491][n491];
        end
    endgenerate
    generate 
        localparam integer d492 = 16;
        for (n492 = 0; n492 < 16; n492 = n492 + 1) 
        begin: outbit492
            assign data_11[n492 + d492*16 + c17*28*16] = data_11_array[c17][d492][n492];
        end
    endgenerate
    generate 
        localparam integer d493 = 17;
        for (n493 = 0; n493 < 16; n493 = n493 + 1) 
        begin: outbit493
            assign data_11[n493 + d493*16 + c17*28*16] = data_11_array[c17][d493][n493];
        end
    endgenerate
    generate 
        localparam integer d494 = 18;
        for (n494 = 0; n494 < 16; n494 = n494 + 1) 
        begin: outbit494
            assign data_11[n494 + d494*16 + c17*28*16] = data_11_array[c17][d494][n494];
        end
    endgenerate
    generate 
        localparam integer d495 = 19;
        for (n495 = 0; n495 < 16; n495 = n495 + 1) 
        begin: outbit495
            assign data_11[n495 + d495*16 + c17*28*16] = data_11_array[c17][d495][n495];
        end
    endgenerate
    generate 
        localparam integer d496 = 20;
        for (n496 = 0; n496 < 16; n496 = n496 + 1) 
        begin: outbit496
            assign data_11[n496 + d496*16 + c17*28*16] = data_11_array[c17][d496][n496];
        end
    endgenerate
    generate 
        localparam integer d497 = 21;
        for (n497 = 0; n497 < 16; n497 = n497 + 1) 
        begin: outbit497
            assign data_11[n497 + d497*16 + c17*28*16] = data_11_array[c17][d497][n497];
        end
    endgenerate
    generate 
        localparam integer d498 = 22;
        for (n498 = 0; n498 < 16; n498 = n498 + 1) 
        begin: outbit498
            assign data_11[n498 + d498*16 + c17*28*16] = data_11_array[c17][d498][n498];
        end
    endgenerate
    generate 
        localparam integer d499 = 23;
        for (n499 = 0; n499 < 16; n499 = n499 + 1) 
        begin: outbit499
            assign data_11[n499 + d499*16 + c17*28*16] = data_11_array[c17][d499][n499];
        end
    endgenerate
    generate 
        localparam integer d500 = 24;
        for (n500 = 0; n500 < 16; n500 = n500 + 1) 
        begin: outbit500
            assign data_11[n500 + d500*16 + c17*28*16] = data_11_array[c17][d500][n500];
        end
    endgenerate
    generate 
        localparam integer d501 = 25;
        for (n501 = 0; n501 < 16; n501 = n501 + 1) 
        begin: outbit501
            assign data_11[n501 + d501*16 + c17*28*16] = data_11_array[c17][d501][n501];
        end
    endgenerate
    generate 
        localparam integer d502 = 26;
        for (n502 = 0; n502 < 16; n502 = n502 + 1) 
        begin: outbit502
            assign data_11[n502 + d502*16 + c17*28*16] = data_11_array[c17][d502][n502];
        end
    endgenerate
    generate 
        localparam integer d503 = 27;
        for (n503 = 0; n503 < 16; n503 = n503 + 1) 
        begin: outbit503
            assign data_11[n503 + d503*16 + c17*28*16] = data_11_array[c17][d503][n503];
        end
    endgenerate
    localparam integer c18 = 18;
    generate 
        localparam integer d504 = 0;
        for (n504 = 0; n504 < 16; n504 = n504 + 1) 
        begin: outbit504
            assign data_11[n504 + d504*16 + c18*28*16] = data_11_array[c18][d504][n504];
        end
    endgenerate
    generate 
        localparam integer d505 = 1;
        for (n505 = 0; n505 < 16; n505 = n505 + 1) 
        begin: outbit505
            assign data_11[n505 + d505*16 + c18*28*16] = data_11_array[c18][d505][n505];
        end
    endgenerate
    generate 
        localparam integer d506 = 2;
        for (n506 = 0; n506 < 16; n506 = n506 + 1) 
        begin: outbit506
            assign data_11[n506 + d506*16 + c18*28*16] = data_11_array[c18][d506][n506];
        end
    endgenerate
    generate 
        localparam integer d507 = 3;
        for (n507 = 0; n507 < 16; n507 = n507 + 1) 
        begin: outbit507
            assign data_11[n507 + d507*16 + c18*28*16] = data_11_array[c18][d507][n507];
        end
    endgenerate
    generate 
        localparam integer d508 = 4;
        for (n508 = 0; n508 < 16; n508 = n508 + 1) 
        begin: outbit508
            assign data_11[n508 + d508*16 + c18*28*16] = data_11_array[c18][d508][n508];
        end
    endgenerate
    generate 
        localparam integer d509 = 5;
        for (n509 = 0; n509 < 16; n509 = n509 + 1) 
        begin: outbit509
            assign data_11[n509 + d509*16 + c18*28*16] = data_11_array[c18][d509][n509];
        end
    endgenerate
    generate 
        localparam integer d510 = 6;
        for (n510 = 0; n510 < 16; n510 = n510 + 1) 
        begin: outbit510
            assign data_11[n510 + d510*16 + c18*28*16] = data_11_array[c18][d510][n510];
        end
    endgenerate
    generate 
        localparam integer d511 = 7;
        for (n511 = 0; n511 < 16; n511 = n511 + 1) 
        begin: outbit511
            assign data_11[n511 + d511*16 + c18*28*16] = data_11_array[c18][d511][n511];
        end
    endgenerate
    generate 
        localparam integer d512 = 8;
        for (n512 = 0; n512 < 16; n512 = n512 + 1) 
        begin: outbit512
            assign data_11[n512 + d512*16 + c18*28*16] = data_11_array[c18][d512][n512];
        end
    endgenerate
    generate 
        localparam integer d513 = 9;
        for (n513 = 0; n513 < 16; n513 = n513 + 1) 
        begin: outbit513
            assign data_11[n513 + d513*16 + c18*28*16] = data_11_array[c18][d513][n513];
        end
    endgenerate
    generate 
        localparam integer d514 = 10;
        for (n514 = 0; n514 < 16; n514 = n514 + 1) 
        begin: outbit514
            assign data_11[n514 + d514*16 + c18*28*16] = data_11_array[c18][d514][n514];
        end
    endgenerate
    generate 
        localparam integer d515 = 11;
        for (n515 = 0; n515 < 16; n515 = n515 + 1) 
        begin: outbit515
            assign data_11[n515 + d515*16 + c18*28*16] = data_11_array[c18][d515][n515];
        end
    endgenerate
    generate 
        localparam integer d516 = 12;
        for (n516 = 0; n516 < 16; n516 = n516 + 1) 
        begin: outbit516
            assign data_11[n516 + d516*16 + c18*28*16] = data_11_array[c18][d516][n516];
        end
    endgenerate
    generate 
        localparam integer d517 = 13;
        for (n517 = 0; n517 < 16; n517 = n517 + 1) 
        begin: outbit517
            assign data_11[n517 + d517*16 + c18*28*16] = data_11_array[c18][d517][n517];
        end
    endgenerate
    generate 
        localparam integer d518 = 14;
        for (n518 = 0; n518 < 16; n518 = n518 + 1) 
        begin: outbit518
            assign data_11[n518 + d518*16 + c18*28*16] = data_11_array[c18][d518][n518];
        end
    endgenerate
    generate 
        localparam integer d519 = 15;
        for (n519 = 0; n519 < 16; n519 = n519 + 1) 
        begin: outbit519
            assign data_11[n519 + d519*16 + c18*28*16] = data_11_array[c18][d519][n519];
        end
    endgenerate
    generate 
        localparam integer d520 = 16;
        for (n520 = 0; n520 < 16; n520 = n520 + 1) 
        begin: outbit520
            assign data_11[n520 + d520*16 + c18*28*16] = data_11_array[c18][d520][n520];
        end
    endgenerate
    generate 
        localparam integer d521 = 17;
        for (n521 = 0; n521 < 16; n521 = n521 + 1) 
        begin: outbit521
            assign data_11[n521 + d521*16 + c18*28*16] = data_11_array[c18][d521][n521];
        end
    endgenerate
    generate 
        localparam integer d522 = 18;
        for (n522 = 0; n522 < 16; n522 = n522 + 1) 
        begin: outbit522
            assign data_11[n522 + d522*16 + c18*28*16] = data_11_array[c18][d522][n522];
        end
    endgenerate
    generate 
        localparam integer d523 = 19;
        for (n523 = 0; n523 < 16; n523 = n523 + 1) 
        begin: outbit523
            assign data_11[n523 + d523*16 + c18*28*16] = data_11_array[c18][d523][n523];
        end
    endgenerate
    generate 
        localparam integer d524 = 20;
        for (n524 = 0; n524 < 16; n524 = n524 + 1) 
        begin: outbit524
            assign data_11[n524 + d524*16 + c18*28*16] = data_11_array[c18][d524][n524];
        end
    endgenerate
    generate 
        localparam integer d525 = 21;
        for (n525 = 0; n525 < 16; n525 = n525 + 1) 
        begin: outbit525
            assign data_11[n525 + d525*16 + c18*28*16] = data_11_array[c18][d525][n525];
        end
    endgenerate
    generate 
        localparam integer d526 = 22;
        for (n526 = 0; n526 < 16; n526 = n526 + 1) 
        begin: outbit526
            assign data_11[n526 + d526*16 + c18*28*16] = data_11_array[c18][d526][n526];
        end
    endgenerate
    generate 
        localparam integer d527 = 23;
        for (n527 = 0; n527 < 16; n527 = n527 + 1) 
        begin: outbit527
            assign data_11[n527 + d527*16 + c18*28*16] = data_11_array[c18][d527][n527];
        end
    endgenerate
    generate 
        localparam integer d528 = 24;
        for (n528 = 0; n528 < 16; n528 = n528 + 1) 
        begin: outbit528
            assign data_11[n528 + d528*16 + c18*28*16] = data_11_array[c18][d528][n528];
        end
    endgenerate
    generate 
        localparam integer d529 = 25;
        for (n529 = 0; n529 < 16; n529 = n529 + 1) 
        begin: outbit529
            assign data_11[n529 + d529*16 + c18*28*16] = data_11_array[c18][d529][n529];
        end
    endgenerate
    generate 
        localparam integer d530 = 26;
        for (n530 = 0; n530 < 16; n530 = n530 + 1) 
        begin: outbit530
            assign data_11[n530 + d530*16 + c18*28*16] = data_11_array[c18][d530][n530];
        end
    endgenerate
    generate 
        localparam integer d531 = 27;
        for (n531 = 0; n531 < 16; n531 = n531 + 1) 
        begin: outbit531
            assign data_11[n531 + d531*16 + c18*28*16] = data_11_array[c18][d531][n531];
        end
    endgenerate
    localparam integer c19 = 19;
    generate 
        localparam integer d532 = 0;
        for (n532 = 0; n532 < 16; n532 = n532 + 1) 
        begin: outbit532
            assign data_11[n532 + d532*16 + c19*28*16] = data_11_array[c19][d532][n532];
        end
    endgenerate
    generate 
        localparam integer d533 = 1;
        for (n533 = 0; n533 < 16; n533 = n533 + 1) 
        begin: outbit533
            assign data_11[n533 + d533*16 + c19*28*16] = data_11_array[c19][d533][n533];
        end
    endgenerate
    generate 
        localparam integer d534 = 2;
        for (n534 = 0; n534 < 16; n534 = n534 + 1) 
        begin: outbit534
            assign data_11[n534 + d534*16 + c19*28*16] = data_11_array[c19][d534][n534];
        end
    endgenerate
    generate 
        localparam integer d535 = 3;
        for (n535 = 0; n535 < 16; n535 = n535 + 1) 
        begin: outbit535
            assign data_11[n535 + d535*16 + c19*28*16] = data_11_array[c19][d535][n535];
        end
    endgenerate
    generate 
        localparam integer d536 = 4;
        for (n536 = 0; n536 < 16; n536 = n536 + 1) 
        begin: outbit536
            assign data_11[n536 + d536*16 + c19*28*16] = data_11_array[c19][d536][n536];
        end
    endgenerate
    generate 
        localparam integer d537 = 5;
        for (n537 = 0; n537 < 16; n537 = n537 + 1) 
        begin: outbit537
            assign data_11[n537 + d537*16 + c19*28*16] = data_11_array[c19][d537][n537];
        end
    endgenerate
    generate 
        localparam integer d538 = 6;
        for (n538 = 0; n538 < 16; n538 = n538 + 1) 
        begin: outbit538
            assign data_11[n538 + d538*16 + c19*28*16] = data_11_array[c19][d538][n538];
        end
    endgenerate
    generate 
        localparam integer d539 = 7;
        for (n539 = 0; n539 < 16; n539 = n539 + 1) 
        begin: outbit539
            assign data_11[n539 + d539*16 + c19*28*16] = data_11_array[c19][d539][n539];
        end
    endgenerate
    generate 
        localparam integer d540 = 8;
        for (n540 = 0; n540 < 16; n540 = n540 + 1) 
        begin: outbit540
            assign data_11[n540 + d540*16 + c19*28*16] = data_11_array[c19][d540][n540];
        end
    endgenerate
    generate 
        localparam integer d541 = 9;
        for (n541 = 0; n541 < 16; n541 = n541 + 1) 
        begin: outbit541
            assign data_11[n541 + d541*16 + c19*28*16] = data_11_array[c19][d541][n541];
        end
    endgenerate
    generate 
        localparam integer d542 = 10;
        for (n542 = 0; n542 < 16; n542 = n542 + 1) 
        begin: outbit542
            assign data_11[n542 + d542*16 + c19*28*16] = data_11_array[c19][d542][n542];
        end
    endgenerate
    generate 
        localparam integer d543 = 11;
        for (n543 = 0; n543 < 16; n543 = n543 + 1) 
        begin: outbit543
            assign data_11[n543 + d543*16 + c19*28*16] = data_11_array[c19][d543][n543];
        end
    endgenerate
    generate 
        localparam integer d544 = 12;
        for (n544 = 0; n544 < 16; n544 = n544 + 1) 
        begin: outbit544
            assign data_11[n544 + d544*16 + c19*28*16] = data_11_array[c19][d544][n544];
        end
    endgenerate
    generate 
        localparam integer d545 = 13;
        for (n545 = 0; n545 < 16; n545 = n545 + 1) 
        begin: outbit545
            assign data_11[n545 + d545*16 + c19*28*16] = data_11_array[c19][d545][n545];
        end
    endgenerate
    generate 
        localparam integer d546 = 14;
        for (n546 = 0; n546 < 16; n546 = n546 + 1) 
        begin: outbit546
            assign data_11[n546 + d546*16 + c19*28*16] = data_11_array[c19][d546][n546];
        end
    endgenerate
    generate 
        localparam integer d547 = 15;
        for (n547 = 0; n547 < 16; n547 = n547 + 1) 
        begin: outbit547
            assign data_11[n547 + d547*16 + c19*28*16] = data_11_array[c19][d547][n547];
        end
    endgenerate
    generate 
        localparam integer d548 = 16;
        for (n548 = 0; n548 < 16; n548 = n548 + 1) 
        begin: outbit548
            assign data_11[n548 + d548*16 + c19*28*16] = data_11_array[c19][d548][n548];
        end
    endgenerate
    generate 
        localparam integer d549 = 17;
        for (n549 = 0; n549 < 16; n549 = n549 + 1) 
        begin: outbit549
            assign data_11[n549 + d549*16 + c19*28*16] = data_11_array[c19][d549][n549];
        end
    endgenerate
    generate 
        localparam integer d550 = 18;
        for (n550 = 0; n550 < 16; n550 = n550 + 1) 
        begin: outbit550
            assign data_11[n550 + d550*16 + c19*28*16] = data_11_array[c19][d550][n550];
        end
    endgenerate
    generate 
        localparam integer d551 = 19;
        for (n551 = 0; n551 < 16; n551 = n551 + 1) 
        begin: outbit551
            assign data_11[n551 + d551*16 + c19*28*16] = data_11_array[c19][d551][n551];
        end
    endgenerate
    generate 
        localparam integer d552 = 20;
        for (n552 = 0; n552 < 16; n552 = n552 + 1) 
        begin: outbit552
            assign data_11[n552 + d552*16 + c19*28*16] = data_11_array[c19][d552][n552];
        end
    endgenerate
    generate 
        localparam integer d553 = 21;
        for (n553 = 0; n553 < 16; n553 = n553 + 1) 
        begin: outbit553
            assign data_11[n553 + d553*16 + c19*28*16] = data_11_array[c19][d553][n553];
        end
    endgenerate
    generate 
        localparam integer d554 = 22;
        for (n554 = 0; n554 < 16; n554 = n554 + 1) 
        begin: outbit554
            assign data_11[n554 + d554*16 + c19*28*16] = data_11_array[c19][d554][n554];
        end
    endgenerate
    generate 
        localparam integer d555 = 23;
        for (n555 = 0; n555 < 16; n555 = n555 + 1) 
        begin: outbit555
            assign data_11[n555 + d555*16 + c19*28*16] = data_11_array[c19][d555][n555];
        end
    endgenerate
    generate 
        localparam integer d556 = 24;
        for (n556 = 0; n556 < 16; n556 = n556 + 1) 
        begin: outbit556
            assign data_11[n556 + d556*16 + c19*28*16] = data_11_array[c19][d556][n556];
        end
    endgenerate
    generate 
        localparam integer d557 = 25;
        for (n557 = 0; n557 < 16; n557 = n557 + 1) 
        begin: outbit557
            assign data_11[n557 + d557*16 + c19*28*16] = data_11_array[c19][d557][n557];
        end
    endgenerate
    generate 
        localparam integer d558 = 26;
        for (n558 = 0; n558 < 16; n558 = n558 + 1) 
        begin: outbit558
            assign data_11[n558 + d558*16 + c19*28*16] = data_11_array[c19][d558][n558];
        end
    endgenerate
    generate 
        localparam integer d559 = 27;
        for (n559 = 0; n559 < 16; n559 = n559 + 1) 
        begin: outbit559
            assign data_11[n559 + d559*16 + c19*28*16] = data_11_array[c19][d559][n559];
        end
    endgenerate
    localparam integer c20 = 20;
    generate 
        localparam integer d560 = 0;
        for (n560 = 0; n560 < 16; n560 = n560 + 1) 
        begin: outbit560
            assign data_11[n560 + d560*16 + c20*28*16] = data_11_array[c20][d560][n560];
        end
    endgenerate
    generate 
        localparam integer d561 = 1;
        for (n561 = 0; n561 < 16; n561 = n561 + 1) 
        begin: outbit561
            assign data_11[n561 + d561*16 + c20*28*16] = data_11_array[c20][d561][n561];
        end
    endgenerate
    generate 
        localparam integer d562 = 2;
        for (n562 = 0; n562 < 16; n562 = n562 + 1) 
        begin: outbit562
            assign data_11[n562 + d562*16 + c20*28*16] = data_11_array[c20][d562][n562];
        end
    endgenerate
    generate 
        localparam integer d563 = 3;
        for (n563 = 0; n563 < 16; n563 = n563 + 1) 
        begin: outbit563
            assign data_11[n563 + d563*16 + c20*28*16] = data_11_array[c20][d563][n563];
        end
    endgenerate
    generate 
        localparam integer d564 = 4;
        for (n564 = 0; n564 < 16; n564 = n564 + 1) 
        begin: outbit564
            assign data_11[n564 + d564*16 + c20*28*16] = data_11_array[c20][d564][n564];
        end
    endgenerate
    generate 
        localparam integer d565 = 5;
        for (n565 = 0; n565 < 16; n565 = n565 + 1) 
        begin: outbit565
            assign data_11[n565 + d565*16 + c20*28*16] = data_11_array[c20][d565][n565];
        end
    endgenerate
    generate 
        localparam integer d566 = 6;
        for (n566 = 0; n566 < 16; n566 = n566 + 1) 
        begin: outbit566
            assign data_11[n566 + d566*16 + c20*28*16] = data_11_array[c20][d566][n566];
        end
    endgenerate
    generate 
        localparam integer d567 = 7;
        for (n567 = 0; n567 < 16; n567 = n567 + 1) 
        begin: outbit567
            assign data_11[n567 + d567*16 + c20*28*16] = data_11_array[c20][d567][n567];
        end
    endgenerate
    generate 
        localparam integer d568 = 8;
        for (n568 = 0; n568 < 16; n568 = n568 + 1) 
        begin: outbit568
            assign data_11[n568 + d568*16 + c20*28*16] = data_11_array[c20][d568][n568];
        end
    endgenerate
    generate 
        localparam integer d569 = 9;
        for (n569 = 0; n569 < 16; n569 = n569 + 1) 
        begin: outbit569
            assign data_11[n569 + d569*16 + c20*28*16] = data_11_array[c20][d569][n569];
        end
    endgenerate
    generate 
        localparam integer d570 = 10;
        for (n570 = 0; n570 < 16; n570 = n570 + 1) 
        begin: outbit570
            assign data_11[n570 + d570*16 + c20*28*16] = data_11_array[c20][d570][n570];
        end
    endgenerate
    generate 
        localparam integer d571 = 11;
        for (n571 = 0; n571 < 16; n571 = n571 + 1) 
        begin: outbit571
            assign data_11[n571 + d571*16 + c20*28*16] = data_11_array[c20][d571][n571];
        end
    endgenerate
    generate 
        localparam integer d572 = 12;
        for (n572 = 0; n572 < 16; n572 = n572 + 1) 
        begin: outbit572
            assign data_11[n572 + d572*16 + c20*28*16] = data_11_array[c20][d572][n572];
        end
    endgenerate
    generate 
        localparam integer d573 = 13;
        for (n573 = 0; n573 < 16; n573 = n573 + 1) 
        begin: outbit573
            assign data_11[n573 + d573*16 + c20*28*16] = data_11_array[c20][d573][n573];
        end
    endgenerate
    generate 
        localparam integer d574 = 14;
        for (n574 = 0; n574 < 16; n574 = n574 + 1) 
        begin: outbit574
            assign data_11[n574 + d574*16 + c20*28*16] = data_11_array[c20][d574][n574];
        end
    endgenerate
    generate 
        localparam integer d575 = 15;
        for (n575 = 0; n575 < 16; n575 = n575 + 1) 
        begin: outbit575
            assign data_11[n575 + d575*16 + c20*28*16] = data_11_array[c20][d575][n575];
        end
    endgenerate
    generate 
        localparam integer d576 = 16;
        for (n576 = 0; n576 < 16; n576 = n576 + 1) 
        begin: outbit576
            assign data_11[n576 + d576*16 + c20*28*16] = data_11_array[c20][d576][n576];
        end
    endgenerate
    generate 
        localparam integer d577 = 17;
        for (n577 = 0; n577 < 16; n577 = n577 + 1) 
        begin: outbit577
            assign data_11[n577 + d577*16 + c20*28*16] = data_11_array[c20][d577][n577];
        end
    endgenerate
    generate 
        localparam integer d578 = 18;
        for (n578 = 0; n578 < 16; n578 = n578 + 1) 
        begin: outbit578
            assign data_11[n578 + d578*16 + c20*28*16] = data_11_array[c20][d578][n578];
        end
    endgenerate
    generate 
        localparam integer d579 = 19;
        for (n579 = 0; n579 < 16; n579 = n579 + 1) 
        begin: outbit579
            assign data_11[n579 + d579*16 + c20*28*16] = data_11_array[c20][d579][n579];
        end
    endgenerate
    generate 
        localparam integer d580 = 20;
        for (n580 = 0; n580 < 16; n580 = n580 + 1) 
        begin: outbit580
            assign data_11[n580 + d580*16 + c20*28*16] = data_11_array[c20][d580][n580];
        end
    endgenerate
    generate 
        localparam integer d581 = 21;
        for (n581 = 0; n581 < 16; n581 = n581 + 1) 
        begin: outbit581
            assign data_11[n581 + d581*16 + c20*28*16] = data_11_array[c20][d581][n581];
        end
    endgenerate
    generate 
        localparam integer d582 = 22;
        for (n582 = 0; n582 < 16; n582 = n582 + 1) 
        begin: outbit582
            assign data_11[n582 + d582*16 + c20*28*16] = data_11_array[c20][d582][n582];
        end
    endgenerate
    generate 
        localparam integer d583 = 23;
        for (n583 = 0; n583 < 16; n583 = n583 + 1) 
        begin: outbit583
            assign data_11[n583 + d583*16 + c20*28*16] = data_11_array[c20][d583][n583];
        end
    endgenerate
    generate 
        localparam integer d584 = 24;
        for (n584 = 0; n584 < 16; n584 = n584 + 1) 
        begin: outbit584
            assign data_11[n584 + d584*16 + c20*28*16] = data_11_array[c20][d584][n584];
        end
    endgenerate
    generate 
        localparam integer d585 = 25;
        for (n585 = 0; n585 < 16; n585 = n585 + 1) 
        begin: outbit585
            assign data_11[n585 + d585*16 + c20*28*16] = data_11_array[c20][d585][n585];
        end
    endgenerate
    generate 
        localparam integer d586 = 26;
        for (n586 = 0; n586 < 16; n586 = n586 + 1) 
        begin: outbit586
            assign data_11[n586 + d586*16 + c20*28*16] = data_11_array[c20][d586][n586];
        end
    endgenerate
    generate 
        localparam integer d587 = 27;
        for (n587 = 0; n587 < 16; n587 = n587 + 1) 
        begin: outbit587
            assign data_11[n587 + d587*16 + c20*28*16] = data_11_array[c20][d587][n587];
        end
    endgenerate
    localparam integer c21 = 21;
    generate 
        localparam integer d588 = 0;
        for (n588 = 0; n588 < 16; n588 = n588 + 1) 
        begin: outbit588
            assign data_11[n588 + d588*16 + c21*28*16] = data_11_array[c21][d588][n588];
        end
    endgenerate
    generate 
        localparam integer d589 = 1;
        for (n589 = 0; n589 < 16; n589 = n589 + 1) 
        begin: outbit589
            assign data_11[n589 + d589*16 + c21*28*16] = data_11_array[c21][d589][n589];
        end
    endgenerate
    generate 
        localparam integer d590 = 2;
        for (n590 = 0; n590 < 16; n590 = n590 + 1) 
        begin: outbit590
            assign data_11[n590 + d590*16 + c21*28*16] = data_11_array[c21][d590][n590];
        end
    endgenerate
    generate 
        localparam integer d591 = 3;
        for (n591 = 0; n591 < 16; n591 = n591 + 1) 
        begin: outbit591
            assign data_11[n591 + d591*16 + c21*28*16] = data_11_array[c21][d591][n591];
        end
    endgenerate
    generate 
        localparam integer d592 = 4;
        for (n592 = 0; n592 < 16; n592 = n592 + 1) 
        begin: outbit592
            assign data_11[n592 + d592*16 + c21*28*16] = data_11_array[c21][d592][n592];
        end
    endgenerate
    generate 
        localparam integer d593 = 5;
        for (n593 = 0; n593 < 16; n593 = n593 + 1) 
        begin: outbit593
            assign data_11[n593 + d593*16 + c21*28*16] = data_11_array[c21][d593][n593];
        end
    endgenerate
    generate 
        localparam integer d594 = 6;
        for (n594 = 0; n594 < 16; n594 = n594 + 1) 
        begin: outbit594
            assign data_11[n594 + d594*16 + c21*28*16] = data_11_array[c21][d594][n594];
        end
    endgenerate
    generate 
        localparam integer d595 = 7;
        for (n595 = 0; n595 < 16; n595 = n595 + 1) 
        begin: outbit595
            assign data_11[n595 + d595*16 + c21*28*16] = data_11_array[c21][d595][n595];
        end
    endgenerate
    generate 
        localparam integer d596 = 8;
        for (n596 = 0; n596 < 16; n596 = n596 + 1) 
        begin: outbit596
            assign data_11[n596 + d596*16 + c21*28*16] = data_11_array[c21][d596][n596];
        end
    endgenerate
    generate 
        localparam integer d597 = 9;
        for (n597 = 0; n597 < 16; n597 = n597 + 1) 
        begin: outbit597
            assign data_11[n597 + d597*16 + c21*28*16] = data_11_array[c21][d597][n597];
        end
    endgenerate
    generate 
        localparam integer d598 = 10;
        for (n598 = 0; n598 < 16; n598 = n598 + 1) 
        begin: outbit598
            assign data_11[n598 + d598*16 + c21*28*16] = data_11_array[c21][d598][n598];
        end
    endgenerate
    generate 
        localparam integer d599 = 11;
        for (n599 = 0; n599 < 16; n599 = n599 + 1) 
        begin: outbit599
            assign data_11[n599 + d599*16 + c21*28*16] = data_11_array[c21][d599][n599];
        end
    endgenerate
    generate 
        localparam integer d600 = 12;
        for (n600 = 0; n600 < 16; n600 = n600 + 1) 
        begin: outbit600
            assign data_11[n600 + d600*16 + c21*28*16] = data_11_array[c21][d600][n600];
        end
    endgenerate
    generate 
        localparam integer d601 = 13;
        for (n601 = 0; n601 < 16; n601 = n601 + 1) 
        begin: outbit601
            assign data_11[n601 + d601*16 + c21*28*16] = data_11_array[c21][d601][n601];
        end
    endgenerate
    generate 
        localparam integer d602 = 14;
        for (n602 = 0; n602 < 16; n602 = n602 + 1) 
        begin: outbit602
            assign data_11[n602 + d602*16 + c21*28*16] = data_11_array[c21][d602][n602];
        end
    endgenerate
    generate 
        localparam integer d603 = 15;
        for (n603 = 0; n603 < 16; n603 = n603 + 1) 
        begin: outbit603
            assign data_11[n603 + d603*16 + c21*28*16] = data_11_array[c21][d603][n603];
        end
    endgenerate
    generate 
        localparam integer d604 = 16;
        for (n604 = 0; n604 < 16; n604 = n604 + 1) 
        begin: outbit604
            assign data_11[n604 + d604*16 + c21*28*16] = data_11_array[c21][d604][n604];
        end
    endgenerate
    generate 
        localparam integer d605 = 17;
        for (n605 = 0; n605 < 16; n605 = n605 + 1) 
        begin: outbit605
            assign data_11[n605 + d605*16 + c21*28*16] = data_11_array[c21][d605][n605];
        end
    endgenerate
    generate 
        localparam integer d606 = 18;
        for (n606 = 0; n606 < 16; n606 = n606 + 1) 
        begin: outbit606
            assign data_11[n606 + d606*16 + c21*28*16] = data_11_array[c21][d606][n606];
        end
    endgenerate
    generate 
        localparam integer d607 = 19;
        for (n607 = 0; n607 < 16; n607 = n607 + 1) 
        begin: outbit607
            assign data_11[n607 + d607*16 + c21*28*16] = data_11_array[c21][d607][n607];
        end
    endgenerate
    generate 
        localparam integer d608 = 20;
        for (n608 = 0; n608 < 16; n608 = n608 + 1) 
        begin: outbit608
            assign data_11[n608 + d608*16 + c21*28*16] = data_11_array[c21][d608][n608];
        end
    endgenerate
    generate 
        localparam integer d609 = 21;
        for (n609 = 0; n609 < 16; n609 = n609 + 1) 
        begin: outbit609
            assign data_11[n609 + d609*16 + c21*28*16] = data_11_array[c21][d609][n609];
        end
    endgenerate
    generate 
        localparam integer d610 = 22;
        for (n610 = 0; n610 < 16; n610 = n610 + 1) 
        begin: outbit610
            assign data_11[n610 + d610*16 + c21*28*16] = data_11_array[c21][d610][n610];
        end
    endgenerate
    generate 
        localparam integer d611 = 23;
        for (n611 = 0; n611 < 16; n611 = n611 + 1) 
        begin: outbit611
            assign data_11[n611 + d611*16 + c21*28*16] = data_11_array[c21][d611][n611];
        end
    endgenerate
    generate 
        localparam integer d612 = 24;
        for (n612 = 0; n612 < 16; n612 = n612 + 1) 
        begin: outbit612
            assign data_11[n612 + d612*16 + c21*28*16] = data_11_array[c21][d612][n612];
        end
    endgenerate
    generate 
        localparam integer d613 = 25;
        for (n613 = 0; n613 < 16; n613 = n613 + 1) 
        begin: outbit613
            assign data_11[n613 + d613*16 + c21*28*16] = data_11_array[c21][d613][n613];
        end
    endgenerate
    generate 
        localparam integer d614 = 26;
        for (n614 = 0; n614 < 16; n614 = n614 + 1) 
        begin: outbit614
            assign data_11[n614 + d614*16 + c21*28*16] = data_11_array[c21][d614][n614];
        end
    endgenerate
    generate 
        localparam integer d615 = 27;
        for (n615 = 0; n615 < 16; n615 = n615 + 1) 
        begin: outbit615
            assign data_11[n615 + d615*16 + c21*28*16] = data_11_array[c21][d615][n615];
        end
    endgenerate
    localparam integer c22 = 22;
    generate 
        localparam integer d616 = 0;
        for (n616 = 0; n616 < 16; n616 = n616 + 1) 
        begin: outbit616
            assign data_11[n616 + d616*16 + c22*28*16] = data_11_array[c22][d616][n616];
        end
    endgenerate
    generate 
        localparam integer d617 = 1;
        for (n617 = 0; n617 < 16; n617 = n617 + 1) 
        begin: outbit617
            assign data_11[n617 + d617*16 + c22*28*16] = data_11_array[c22][d617][n617];
        end
    endgenerate
    generate 
        localparam integer d618 = 2;
        for (n618 = 0; n618 < 16; n618 = n618 + 1) 
        begin: outbit618
            assign data_11[n618 + d618*16 + c22*28*16] = data_11_array[c22][d618][n618];
        end
    endgenerate
    generate 
        localparam integer d619 = 3;
        for (n619 = 0; n619 < 16; n619 = n619 + 1) 
        begin: outbit619
            assign data_11[n619 + d619*16 + c22*28*16] = data_11_array[c22][d619][n619];
        end
    endgenerate
    generate 
        localparam integer d620 = 4;
        for (n620 = 0; n620 < 16; n620 = n620 + 1) 
        begin: outbit620
            assign data_11[n620 + d620*16 + c22*28*16] = data_11_array[c22][d620][n620];
        end
    endgenerate
    generate 
        localparam integer d621 = 5;
        for (n621 = 0; n621 < 16; n621 = n621 + 1) 
        begin: outbit621
            assign data_11[n621 + d621*16 + c22*28*16] = data_11_array[c22][d621][n621];
        end
    endgenerate
    generate 
        localparam integer d622 = 6;
        for (n622 = 0; n622 < 16; n622 = n622 + 1) 
        begin: outbit622
            assign data_11[n622 + d622*16 + c22*28*16] = data_11_array[c22][d622][n622];
        end
    endgenerate
    generate 
        localparam integer d623 = 7;
        for (n623 = 0; n623 < 16; n623 = n623 + 1) 
        begin: outbit623
            assign data_11[n623 + d623*16 + c22*28*16] = data_11_array[c22][d623][n623];
        end
    endgenerate
    generate 
        localparam integer d624 = 8;
        for (n624 = 0; n624 < 16; n624 = n624 + 1) 
        begin: outbit624
            assign data_11[n624 + d624*16 + c22*28*16] = data_11_array[c22][d624][n624];
        end
    endgenerate
    generate 
        localparam integer d625 = 9;
        for (n625 = 0; n625 < 16; n625 = n625 + 1) 
        begin: outbit625
            assign data_11[n625 + d625*16 + c22*28*16] = data_11_array[c22][d625][n625];
        end
    endgenerate
    generate 
        localparam integer d626 = 10;
        for (n626 = 0; n626 < 16; n626 = n626 + 1) 
        begin: outbit626
            assign data_11[n626 + d626*16 + c22*28*16] = data_11_array[c22][d626][n626];
        end
    endgenerate
    generate 
        localparam integer d627 = 11;
        for (n627 = 0; n627 < 16; n627 = n627 + 1) 
        begin: outbit627
            assign data_11[n627 + d627*16 + c22*28*16] = data_11_array[c22][d627][n627];
        end
    endgenerate
    generate 
        localparam integer d628 = 12;
        for (n628 = 0; n628 < 16; n628 = n628 + 1) 
        begin: outbit628
            assign data_11[n628 + d628*16 + c22*28*16] = data_11_array[c22][d628][n628];
        end
    endgenerate
    generate 
        localparam integer d629 = 13;
        for (n629 = 0; n629 < 16; n629 = n629 + 1) 
        begin: outbit629
            assign data_11[n629 + d629*16 + c22*28*16] = data_11_array[c22][d629][n629];
        end
    endgenerate
    generate 
        localparam integer d630 = 14;
        for (n630 = 0; n630 < 16; n630 = n630 + 1) 
        begin: outbit630
            assign data_11[n630 + d630*16 + c22*28*16] = data_11_array[c22][d630][n630];
        end
    endgenerate
    generate 
        localparam integer d631 = 15;
        for (n631 = 0; n631 < 16; n631 = n631 + 1) 
        begin: outbit631
            assign data_11[n631 + d631*16 + c22*28*16] = data_11_array[c22][d631][n631];
        end
    endgenerate
    generate 
        localparam integer d632 = 16;
        for (n632 = 0; n632 < 16; n632 = n632 + 1) 
        begin: outbit632
            assign data_11[n632 + d632*16 + c22*28*16] = data_11_array[c22][d632][n632];
        end
    endgenerate
    generate 
        localparam integer d633 = 17;
        for (n633 = 0; n633 < 16; n633 = n633 + 1) 
        begin: outbit633
            assign data_11[n633 + d633*16 + c22*28*16] = data_11_array[c22][d633][n633];
        end
    endgenerate
    generate 
        localparam integer d634 = 18;
        for (n634 = 0; n634 < 16; n634 = n634 + 1) 
        begin: outbit634
            assign data_11[n634 + d634*16 + c22*28*16] = data_11_array[c22][d634][n634];
        end
    endgenerate
    generate 
        localparam integer d635 = 19;
        for (n635 = 0; n635 < 16; n635 = n635 + 1) 
        begin: outbit635
            assign data_11[n635 + d635*16 + c22*28*16] = data_11_array[c22][d635][n635];
        end
    endgenerate
    generate 
        localparam integer d636 = 20;
        for (n636 = 0; n636 < 16; n636 = n636 + 1) 
        begin: outbit636
            assign data_11[n636 + d636*16 + c22*28*16] = data_11_array[c22][d636][n636];
        end
    endgenerate
    generate 
        localparam integer d637 = 21;
        for (n637 = 0; n637 < 16; n637 = n637 + 1) 
        begin: outbit637
            assign data_11[n637 + d637*16 + c22*28*16] = data_11_array[c22][d637][n637];
        end
    endgenerate
    generate 
        localparam integer d638 = 22;
        for (n638 = 0; n638 < 16; n638 = n638 + 1) 
        begin: outbit638
            assign data_11[n638 + d638*16 + c22*28*16] = data_11_array[c22][d638][n638];
        end
    endgenerate
    generate 
        localparam integer d639 = 23;
        for (n639 = 0; n639 < 16; n639 = n639 + 1) 
        begin: outbit639
            assign data_11[n639 + d639*16 + c22*28*16] = data_11_array[c22][d639][n639];
        end
    endgenerate
    generate 
        localparam integer d640 = 24;
        for (n640 = 0; n640 < 16; n640 = n640 + 1) 
        begin: outbit640
            assign data_11[n640 + d640*16 + c22*28*16] = data_11_array[c22][d640][n640];
        end
    endgenerate
    generate 
        localparam integer d641 = 25;
        for (n641 = 0; n641 < 16; n641 = n641 + 1) 
        begin: outbit641
            assign data_11[n641 + d641*16 + c22*28*16] = data_11_array[c22][d641][n641];
        end
    endgenerate
    generate 
        localparam integer d642 = 26;
        for (n642 = 0; n642 < 16; n642 = n642 + 1) 
        begin: outbit642
            assign data_11[n642 + d642*16 + c22*28*16] = data_11_array[c22][d642][n642];
        end
    endgenerate
    generate 
        localparam integer d643 = 27;
        for (n643 = 0; n643 < 16; n643 = n643 + 1) 
        begin: outbit643
            assign data_11[n643 + d643*16 + c22*28*16] = data_11_array[c22][d643][n643];
        end
    endgenerate
    localparam integer c23 = 23;
    generate 
        localparam integer d644 = 0;
        for (n644 = 0; n644 < 16; n644 = n644 + 1) 
        begin: outbit644
            assign data_11[n644 + d644*16 + c23*28*16] = data_11_array[c23][d644][n644];
        end
    endgenerate
    generate 
        localparam integer d645 = 1;
        for (n645 = 0; n645 < 16; n645 = n645 + 1) 
        begin: outbit645
            assign data_11[n645 + d645*16 + c23*28*16] = data_11_array[c23][d645][n645];
        end
    endgenerate
    generate 
        localparam integer d646 = 2;
        for (n646 = 0; n646 < 16; n646 = n646 + 1) 
        begin: outbit646
            assign data_11[n646 + d646*16 + c23*28*16] = data_11_array[c23][d646][n646];
        end
    endgenerate
    generate 
        localparam integer d647 = 3;
        for (n647 = 0; n647 < 16; n647 = n647 + 1) 
        begin: outbit647
            assign data_11[n647 + d647*16 + c23*28*16] = data_11_array[c23][d647][n647];
        end
    endgenerate
    generate 
        localparam integer d648 = 4;
        for (n648 = 0; n648 < 16; n648 = n648 + 1) 
        begin: outbit648
            assign data_11[n648 + d648*16 + c23*28*16] = data_11_array[c23][d648][n648];
        end
    endgenerate
    generate 
        localparam integer d649 = 5;
        for (n649 = 0; n649 < 16; n649 = n649 + 1) 
        begin: outbit649
            assign data_11[n649 + d649*16 + c23*28*16] = data_11_array[c23][d649][n649];
        end
    endgenerate
    generate 
        localparam integer d650 = 6;
        for (n650 = 0; n650 < 16; n650 = n650 + 1) 
        begin: outbit650
            assign data_11[n650 + d650*16 + c23*28*16] = data_11_array[c23][d650][n650];
        end
    endgenerate
    generate 
        localparam integer d651 = 7;
        for (n651 = 0; n651 < 16; n651 = n651 + 1) 
        begin: outbit651
            assign data_11[n651 + d651*16 + c23*28*16] = data_11_array[c23][d651][n651];
        end
    endgenerate
    generate 
        localparam integer d652 = 8;
        for (n652 = 0; n652 < 16; n652 = n652 + 1) 
        begin: outbit652
            assign data_11[n652 + d652*16 + c23*28*16] = data_11_array[c23][d652][n652];
        end
    endgenerate
    generate 
        localparam integer d653 = 9;
        for (n653 = 0; n653 < 16; n653 = n653 + 1) 
        begin: outbit653
            assign data_11[n653 + d653*16 + c23*28*16] = data_11_array[c23][d653][n653];
        end
    endgenerate
    generate 
        localparam integer d654 = 10;
        for (n654 = 0; n654 < 16; n654 = n654 + 1) 
        begin: outbit654
            assign data_11[n654 + d654*16 + c23*28*16] = data_11_array[c23][d654][n654];
        end
    endgenerate
    generate 
        localparam integer d655 = 11;
        for (n655 = 0; n655 < 16; n655 = n655 + 1) 
        begin: outbit655
            assign data_11[n655 + d655*16 + c23*28*16] = data_11_array[c23][d655][n655];
        end
    endgenerate
    generate 
        localparam integer d656 = 12;
        for (n656 = 0; n656 < 16; n656 = n656 + 1) 
        begin: outbit656
            assign data_11[n656 + d656*16 + c23*28*16] = data_11_array[c23][d656][n656];
        end
    endgenerate
    generate 
        localparam integer d657 = 13;
        for (n657 = 0; n657 < 16; n657 = n657 + 1) 
        begin: outbit657
            assign data_11[n657 + d657*16 + c23*28*16] = data_11_array[c23][d657][n657];
        end
    endgenerate
    generate 
        localparam integer d658 = 14;
        for (n658 = 0; n658 < 16; n658 = n658 + 1) 
        begin: outbit658
            assign data_11[n658 + d658*16 + c23*28*16] = data_11_array[c23][d658][n658];
        end
    endgenerate
    generate 
        localparam integer d659 = 15;
        for (n659 = 0; n659 < 16; n659 = n659 + 1) 
        begin: outbit659
            assign data_11[n659 + d659*16 + c23*28*16] = data_11_array[c23][d659][n659];
        end
    endgenerate
    generate 
        localparam integer d660 = 16;
        for (n660 = 0; n660 < 16; n660 = n660 + 1) 
        begin: outbit660
            assign data_11[n660 + d660*16 + c23*28*16] = data_11_array[c23][d660][n660];
        end
    endgenerate
    generate 
        localparam integer d661 = 17;
        for (n661 = 0; n661 < 16; n661 = n661 + 1) 
        begin: outbit661
            assign data_11[n661 + d661*16 + c23*28*16] = data_11_array[c23][d661][n661];
        end
    endgenerate
    generate 
        localparam integer d662 = 18;
        for (n662 = 0; n662 < 16; n662 = n662 + 1) 
        begin: outbit662
            assign data_11[n662 + d662*16 + c23*28*16] = data_11_array[c23][d662][n662];
        end
    endgenerate
    generate 
        localparam integer d663 = 19;
        for (n663 = 0; n663 < 16; n663 = n663 + 1) 
        begin: outbit663
            assign data_11[n663 + d663*16 + c23*28*16] = data_11_array[c23][d663][n663];
        end
    endgenerate
    generate 
        localparam integer d664 = 20;
        for (n664 = 0; n664 < 16; n664 = n664 + 1) 
        begin: outbit664
            assign data_11[n664 + d664*16 + c23*28*16] = data_11_array[c23][d664][n664];
        end
    endgenerate
    generate 
        localparam integer d665 = 21;
        for (n665 = 0; n665 < 16; n665 = n665 + 1) 
        begin: outbit665
            assign data_11[n665 + d665*16 + c23*28*16] = data_11_array[c23][d665][n665];
        end
    endgenerate
    generate 
        localparam integer d666 = 22;
        for (n666 = 0; n666 < 16; n666 = n666 + 1) 
        begin: outbit666
            assign data_11[n666 + d666*16 + c23*28*16] = data_11_array[c23][d666][n666];
        end
    endgenerate
    generate 
        localparam integer d667 = 23;
        for (n667 = 0; n667 < 16; n667 = n667 + 1) 
        begin: outbit667
            assign data_11[n667 + d667*16 + c23*28*16] = data_11_array[c23][d667][n667];
        end
    endgenerate
    generate 
        localparam integer d668 = 24;
        for (n668 = 0; n668 < 16; n668 = n668 + 1) 
        begin: outbit668
            assign data_11[n668 + d668*16 + c23*28*16] = data_11_array[c23][d668][n668];
        end
    endgenerate
    generate 
        localparam integer d669 = 25;
        for (n669 = 0; n669 < 16; n669 = n669 + 1) 
        begin: outbit669
            assign data_11[n669 + d669*16 + c23*28*16] = data_11_array[c23][d669][n669];
        end
    endgenerate
    generate 
        localparam integer d670 = 26;
        for (n670 = 0; n670 < 16; n670 = n670 + 1) 
        begin: outbit670
            assign data_11[n670 + d670*16 + c23*28*16] = data_11_array[c23][d670][n670];
        end
    endgenerate
    generate 
        localparam integer d671 = 27;
        for (n671 = 0; n671 < 16; n671 = n671 + 1) 
        begin: outbit671
            assign data_11[n671 + d671*16 + c23*28*16] = data_11_array[c23][d671][n671];
        end
    endgenerate
    localparam integer c24 = 24;
    generate 
        localparam integer d672 = 0;
        for (n672 = 0; n672 < 16; n672 = n672 + 1) 
        begin: outbit672
            assign data_11[n672 + d672*16 + c24*28*16] = data_11_array[c24][d672][n672];
        end
    endgenerate
    generate 
        localparam integer d673 = 1;
        for (n673 = 0; n673 < 16; n673 = n673 + 1) 
        begin: outbit673
            assign data_11[n673 + d673*16 + c24*28*16] = data_11_array[c24][d673][n673];
        end
    endgenerate
    generate 
        localparam integer d674 = 2;
        for (n674 = 0; n674 < 16; n674 = n674 + 1) 
        begin: outbit674
            assign data_11[n674 + d674*16 + c24*28*16] = data_11_array[c24][d674][n674];
        end
    endgenerate
    generate 
        localparam integer d675 = 3;
        for (n675 = 0; n675 < 16; n675 = n675 + 1) 
        begin: outbit675
            assign data_11[n675 + d675*16 + c24*28*16] = data_11_array[c24][d675][n675];
        end
    endgenerate
    generate 
        localparam integer d676 = 4;
        for (n676 = 0; n676 < 16; n676 = n676 + 1) 
        begin: outbit676
            assign data_11[n676 + d676*16 + c24*28*16] = data_11_array[c24][d676][n676];
        end
    endgenerate
    generate 
        localparam integer d677 = 5;
        for (n677 = 0; n677 < 16; n677 = n677 + 1) 
        begin: outbit677
            assign data_11[n677 + d677*16 + c24*28*16] = data_11_array[c24][d677][n677];
        end
    endgenerate
    generate 
        localparam integer d678 = 6;
        for (n678 = 0; n678 < 16; n678 = n678 + 1) 
        begin: outbit678
            assign data_11[n678 + d678*16 + c24*28*16] = data_11_array[c24][d678][n678];
        end
    endgenerate
    generate 
        localparam integer d679 = 7;
        for (n679 = 0; n679 < 16; n679 = n679 + 1) 
        begin: outbit679
            assign data_11[n679 + d679*16 + c24*28*16] = data_11_array[c24][d679][n679];
        end
    endgenerate
    generate 
        localparam integer d680 = 8;
        for (n680 = 0; n680 < 16; n680 = n680 + 1) 
        begin: outbit680
            assign data_11[n680 + d680*16 + c24*28*16] = data_11_array[c24][d680][n680];
        end
    endgenerate
    generate 
        localparam integer d681 = 9;
        for (n681 = 0; n681 < 16; n681 = n681 + 1) 
        begin: outbit681
            assign data_11[n681 + d681*16 + c24*28*16] = data_11_array[c24][d681][n681];
        end
    endgenerate
    generate 
        localparam integer d682 = 10;
        for (n682 = 0; n682 < 16; n682 = n682 + 1) 
        begin: outbit682
            assign data_11[n682 + d682*16 + c24*28*16] = data_11_array[c24][d682][n682];
        end
    endgenerate
    generate 
        localparam integer d683 = 11;
        for (n683 = 0; n683 < 16; n683 = n683 + 1) 
        begin: outbit683
            assign data_11[n683 + d683*16 + c24*28*16] = data_11_array[c24][d683][n683];
        end
    endgenerate
    generate 
        localparam integer d684 = 12;
        for (n684 = 0; n684 < 16; n684 = n684 + 1) 
        begin: outbit684
            assign data_11[n684 + d684*16 + c24*28*16] = data_11_array[c24][d684][n684];
        end
    endgenerate
    generate 
        localparam integer d685 = 13;
        for (n685 = 0; n685 < 16; n685 = n685 + 1) 
        begin: outbit685
            assign data_11[n685 + d685*16 + c24*28*16] = data_11_array[c24][d685][n685];
        end
    endgenerate
    generate 
        localparam integer d686 = 14;
        for (n686 = 0; n686 < 16; n686 = n686 + 1) 
        begin: outbit686
            assign data_11[n686 + d686*16 + c24*28*16] = data_11_array[c24][d686][n686];
        end
    endgenerate
    generate 
        localparam integer d687 = 15;
        for (n687 = 0; n687 < 16; n687 = n687 + 1) 
        begin: outbit687
            assign data_11[n687 + d687*16 + c24*28*16] = data_11_array[c24][d687][n687];
        end
    endgenerate
    generate 
        localparam integer d688 = 16;
        for (n688 = 0; n688 < 16; n688 = n688 + 1) 
        begin: outbit688
            assign data_11[n688 + d688*16 + c24*28*16] = data_11_array[c24][d688][n688];
        end
    endgenerate
    generate 
        localparam integer d689 = 17;
        for (n689 = 0; n689 < 16; n689 = n689 + 1) 
        begin: outbit689
            assign data_11[n689 + d689*16 + c24*28*16] = data_11_array[c24][d689][n689];
        end
    endgenerate
    generate 
        localparam integer d690 = 18;
        for (n690 = 0; n690 < 16; n690 = n690 + 1) 
        begin: outbit690
            assign data_11[n690 + d690*16 + c24*28*16] = data_11_array[c24][d690][n690];
        end
    endgenerate
    generate 
        localparam integer d691 = 19;
        for (n691 = 0; n691 < 16; n691 = n691 + 1) 
        begin: outbit691
            assign data_11[n691 + d691*16 + c24*28*16] = data_11_array[c24][d691][n691];
        end
    endgenerate
    generate 
        localparam integer d692 = 20;
        for (n692 = 0; n692 < 16; n692 = n692 + 1) 
        begin: outbit692
            assign data_11[n692 + d692*16 + c24*28*16] = data_11_array[c24][d692][n692];
        end
    endgenerate
    generate 
        localparam integer d693 = 21;
        for (n693 = 0; n693 < 16; n693 = n693 + 1) 
        begin: outbit693
            assign data_11[n693 + d693*16 + c24*28*16] = data_11_array[c24][d693][n693];
        end
    endgenerate
    generate 
        localparam integer d694 = 22;
        for (n694 = 0; n694 < 16; n694 = n694 + 1) 
        begin: outbit694
            assign data_11[n694 + d694*16 + c24*28*16] = data_11_array[c24][d694][n694];
        end
    endgenerate
    generate 
        localparam integer d695 = 23;
        for (n695 = 0; n695 < 16; n695 = n695 + 1) 
        begin: outbit695
            assign data_11[n695 + d695*16 + c24*28*16] = data_11_array[c24][d695][n695];
        end
    endgenerate
    generate 
        localparam integer d696 = 24;
        for (n696 = 0; n696 < 16; n696 = n696 + 1) 
        begin: outbit696
            assign data_11[n696 + d696*16 + c24*28*16] = data_11_array[c24][d696][n696];
        end
    endgenerate
    generate 
        localparam integer d697 = 25;
        for (n697 = 0; n697 < 16; n697 = n697 + 1) 
        begin: outbit697
            assign data_11[n697 + d697*16 + c24*28*16] = data_11_array[c24][d697][n697];
        end
    endgenerate
    generate 
        localparam integer d698 = 26;
        for (n698 = 0; n698 < 16; n698 = n698 + 1) 
        begin: outbit698
            assign data_11[n698 + d698*16 + c24*28*16] = data_11_array[c24][d698][n698];
        end
    endgenerate
    generate 
        localparam integer d699 = 27;
        for (n699 = 0; n699 < 16; n699 = n699 + 1) 
        begin: outbit699
            assign data_11[n699 + d699*16 + c24*28*16] = data_11_array[c24][d699][n699];
        end
    endgenerate
    localparam integer c25 = 25;
    generate 
        localparam integer d700 = 0;
        for (n700 = 0; n700 < 16; n700 = n700 + 1) 
        begin: outbit700
            assign data_11[n700 + d700*16 + c25*28*16] = data_11_array[c25][d700][n700];
        end
    endgenerate
    generate 
        localparam integer d701 = 1;
        for (n701 = 0; n701 < 16; n701 = n701 + 1) 
        begin: outbit701
            assign data_11[n701 + d701*16 + c25*28*16] = data_11_array[c25][d701][n701];
        end
    endgenerate
    generate 
        localparam integer d702 = 2;
        for (n702 = 0; n702 < 16; n702 = n702 + 1) 
        begin: outbit702
            assign data_11[n702 + d702*16 + c25*28*16] = data_11_array[c25][d702][n702];
        end
    endgenerate
    generate 
        localparam integer d703 = 3;
        for (n703 = 0; n703 < 16; n703 = n703 + 1) 
        begin: outbit703
            assign data_11[n703 + d703*16 + c25*28*16] = data_11_array[c25][d703][n703];
        end
    endgenerate
    generate 
        localparam integer d704 = 4;
        for (n704 = 0; n704 < 16; n704 = n704 + 1) 
        begin: outbit704
            assign data_11[n704 + d704*16 + c25*28*16] = data_11_array[c25][d704][n704];
        end
    endgenerate
    generate 
        localparam integer d705 = 5;
        for (n705 = 0; n705 < 16; n705 = n705 + 1) 
        begin: outbit705
            assign data_11[n705 + d705*16 + c25*28*16] = data_11_array[c25][d705][n705];
        end
    endgenerate
    generate 
        localparam integer d706 = 6;
        for (n706 = 0; n706 < 16; n706 = n706 + 1) 
        begin: outbit706
            assign data_11[n706 + d706*16 + c25*28*16] = data_11_array[c25][d706][n706];
        end
    endgenerate
    generate 
        localparam integer d707 = 7;
        for (n707 = 0; n707 < 16; n707 = n707 + 1) 
        begin: outbit707
            assign data_11[n707 + d707*16 + c25*28*16] = data_11_array[c25][d707][n707];
        end
    endgenerate
    generate 
        localparam integer d708 = 8;
        for (n708 = 0; n708 < 16; n708 = n708 + 1) 
        begin: outbit708
            assign data_11[n708 + d708*16 + c25*28*16] = data_11_array[c25][d708][n708];
        end
    endgenerate
    generate 
        localparam integer d709 = 9;
        for (n709 = 0; n709 < 16; n709 = n709 + 1) 
        begin: outbit709
            assign data_11[n709 + d709*16 + c25*28*16] = data_11_array[c25][d709][n709];
        end
    endgenerate
    generate 
        localparam integer d710 = 10;
        for (n710 = 0; n710 < 16; n710 = n710 + 1) 
        begin: outbit710
            assign data_11[n710 + d710*16 + c25*28*16] = data_11_array[c25][d710][n710];
        end
    endgenerate
    generate 
        localparam integer d711 = 11;
        for (n711 = 0; n711 < 16; n711 = n711 + 1) 
        begin: outbit711
            assign data_11[n711 + d711*16 + c25*28*16] = data_11_array[c25][d711][n711];
        end
    endgenerate
    generate 
        localparam integer d712 = 12;
        for (n712 = 0; n712 < 16; n712 = n712 + 1) 
        begin: outbit712
            assign data_11[n712 + d712*16 + c25*28*16] = data_11_array[c25][d712][n712];
        end
    endgenerate
    generate 
        localparam integer d713 = 13;
        for (n713 = 0; n713 < 16; n713 = n713 + 1) 
        begin: outbit713
            assign data_11[n713 + d713*16 + c25*28*16] = data_11_array[c25][d713][n713];
        end
    endgenerate
    generate 
        localparam integer d714 = 14;
        for (n714 = 0; n714 < 16; n714 = n714 + 1) 
        begin: outbit714
            assign data_11[n714 + d714*16 + c25*28*16] = data_11_array[c25][d714][n714];
        end
    endgenerate
    generate 
        localparam integer d715 = 15;
        for (n715 = 0; n715 < 16; n715 = n715 + 1) 
        begin: outbit715
            assign data_11[n715 + d715*16 + c25*28*16] = data_11_array[c25][d715][n715];
        end
    endgenerate
    generate 
        localparam integer d716 = 16;
        for (n716 = 0; n716 < 16; n716 = n716 + 1) 
        begin: outbit716
            assign data_11[n716 + d716*16 + c25*28*16] = data_11_array[c25][d716][n716];
        end
    endgenerate
    generate 
        localparam integer d717 = 17;
        for (n717 = 0; n717 < 16; n717 = n717 + 1) 
        begin: outbit717
            assign data_11[n717 + d717*16 + c25*28*16] = data_11_array[c25][d717][n717];
        end
    endgenerate
    generate 
        localparam integer d718 = 18;
        for (n718 = 0; n718 < 16; n718 = n718 + 1) 
        begin: outbit718
            assign data_11[n718 + d718*16 + c25*28*16] = data_11_array[c25][d718][n718];
        end
    endgenerate
    generate 
        localparam integer d719 = 19;
        for (n719 = 0; n719 < 16; n719 = n719 + 1) 
        begin: outbit719
            assign data_11[n719 + d719*16 + c25*28*16] = data_11_array[c25][d719][n719];
        end
    endgenerate
    generate 
        localparam integer d720 = 20;
        for (n720 = 0; n720 < 16; n720 = n720 + 1) 
        begin: outbit720
            assign data_11[n720 + d720*16 + c25*28*16] = data_11_array[c25][d720][n720];
        end
    endgenerate
    generate 
        localparam integer d721 = 21;
        for (n721 = 0; n721 < 16; n721 = n721 + 1) 
        begin: outbit721
            assign data_11[n721 + d721*16 + c25*28*16] = data_11_array[c25][d721][n721];
        end
    endgenerate
    generate 
        localparam integer d722 = 22;
        for (n722 = 0; n722 < 16; n722 = n722 + 1) 
        begin: outbit722
            assign data_11[n722 + d722*16 + c25*28*16] = data_11_array[c25][d722][n722];
        end
    endgenerate
    generate 
        localparam integer d723 = 23;
        for (n723 = 0; n723 < 16; n723 = n723 + 1) 
        begin: outbit723
            assign data_11[n723 + d723*16 + c25*28*16] = data_11_array[c25][d723][n723];
        end
    endgenerate
    generate 
        localparam integer d724 = 24;
        for (n724 = 0; n724 < 16; n724 = n724 + 1) 
        begin: outbit724
            assign data_11[n724 + d724*16 + c25*28*16] = data_11_array[c25][d724][n724];
        end
    endgenerate
    generate 
        localparam integer d725 = 25;
        for (n725 = 0; n725 < 16; n725 = n725 + 1) 
        begin: outbit725
            assign data_11[n725 + d725*16 + c25*28*16] = data_11_array[c25][d725][n725];
        end
    endgenerate
    generate 
        localparam integer d726 = 26;
        for (n726 = 0; n726 < 16; n726 = n726 + 1) 
        begin: outbit726
            assign data_11[n726 + d726*16 + c25*28*16] = data_11_array[c25][d726][n726];
        end
    endgenerate
    generate 
        localparam integer d727 = 27;
        for (n727 = 0; n727 < 16; n727 = n727 + 1) 
        begin: outbit727
            assign data_11[n727 + d727*16 + c25*28*16] = data_11_array[c25][d727][n727];
        end
    endgenerate
    localparam integer c26 = 26;
    generate 
        localparam integer d728 = 0;
        for (n728 = 0; n728 < 16; n728 = n728 + 1) 
        begin: outbit728
            assign data_11[n728 + d728*16 + c26*28*16] = data_11_array[c26][d728][n728];
        end
    endgenerate
    generate 
        localparam integer d729 = 1;
        for (n729 = 0; n729 < 16; n729 = n729 + 1) 
        begin: outbit729
            assign data_11[n729 + d729*16 + c26*28*16] = data_11_array[c26][d729][n729];
        end
    endgenerate
    generate 
        localparam integer d730 = 2;
        for (n730 = 0; n730 < 16; n730 = n730 + 1) 
        begin: outbit730
            assign data_11[n730 + d730*16 + c26*28*16] = data_11_array[c26][d730][n730];
        end
    endgenerate
    generate 
        localparam integer d731 = 3;
        for (n731 = 0; n731 < 16; n731 = n731 + 1) 
        begin: outbit731
            assign data_11[n731 + d731*16 + c26*28*16] = data_11_array[c26][d731][n731];
        end
    endgenerate
    generate 
        localparam integer d732 = 4;
        for (n732 = 0; n732 < 16; n732 = n732 + 1) 
        begin: outbit732
            assign data_11[n732 + d732*16 + c26*28*16] = data_11_array[c26][d732][n732];
        end
    endgenerate
    generate 
        localparam integer d733 = 5;
        for (n733 = 0; n733 < 16; n733 = n733 + 1) 
        begin: outbit733
            assign data_11[n733 + d733*16 + c26*28*16] = data_11_array[c26][d733][n733];
        end
    endgenerate
    generate 
        localparam integer d734 = 6;
        for (n734 = 0; n734 < 16; n734 = n734 + 1) 
        begin: outbit734
            assign data_11[n734 + d734*16 + c26*28*16] = data_11_array[c26][d734][n734];
        end
    endgenerate
    generate 
        localparam integer d735 = 7;
        for (n735 = 0; n735 < 16; n735 = n735 + 1) 
        begin: outbit735
            assign data_11[n735 + d735*16 + c26*28*16] = data_11_array[c26][d735][n735];
        end
    endgenerate
    generate 
        localparam integer d736 = 8;
        for (n736 = 0; n736 < 16; n736 = n736 + 1) 
        begin: outbit736
            assign data_11[n736 + d736*16 + c26*28*16] = data_11_array[c26][d736][n736];
        end
    endgenerate
    generate 
        localparam integer d737 = 9;
        for (n737 = 0; n737 < 16; n737 = n737 + 1) 
        begin: outbit737
            assign data_11[n737 + d737*16 + c26*28*16] = data_11_array[c26][d737][n737];
        end
    endgenerate
    generate 
        localparam integer d738 = 10;
        for (n738 = 0; n738 < 16; n738 = n738 + 1) 
        begin: outbit738
            assign data_11[n738 + d738*16 + c26*28*16] = data_11_array[c26][d738][n738];
        end
    endgenerate
    generate 
        localparam integer d739 = 11;
        for (n739 = 0; n739 < 16; n739 = n739 + 1) 
        begin: outbit739
            assign data_11[n739 + d739*16 + c26*28*16] = data_11_array[c26][d739][n739];
        end
    endgenerate
    generate 
        localparam integer d740 = 12;
        for (n740 = 0; n740 < 16; n740 = n740 + 1) 
        begin: outbit740
            assign data_11[n740 + d740*16 + c26*28*16] = data_11_array[c26][d740][n740];
        end
    endgenerate
    generate 
        localparam integer d741 = 13;
        for (n741 = 0; n741 < 16; n741 = n741 + 1) 
        begin: outbit741
            assign data_11[n741 + d741*16 + c26*28*16] = data_11_array[c26][d741][n741];
        end
    endgenerate
    generate 
        localparam integer d742 = 14;
        for (n742 = 0; n742 < 16; n742 = n742 + 1) 
        begin: outbit742
            assign data_11[n742 + d742*16 + c26*28*16] = data_11_array[c26][d742][n742];
        end
    endgenerate
    generate 
        localparam integer d743 = 15;
        for (n743 = 0; n743 < 16; n743 = n743 + 1) 
        begin: outbit743
            assign data_11[n743 + d743*16 + c26*28*16] = data_11_array[c26][d743][n743];
        end
    endgenerate
    generate 
        localparam integer d744 = 16;
        for (n744 = 0; n744 < 16; n744 = n744 + 1) 
        begin: outbit744
            assign data_11[n744 + d744*16 + c26*28*16] = data_11_array[c26][d744][n744];
        end
    endgenerate
    generate 
        localparam integer d745 = 17;
        for (n745 = 0; n745 < 16; n745 = n745 + 1) 
        begin: outbit745
            assign data_11[n745 + d745*16 + c26*28*16] = data_11_array[c26][d745][n745];
        end
    endgenerate
    generate 
        localparam integer d746 = 18;
        for (n746 = 0; n746 < 16; n746 = n746 + 1) 
        begin: outbit746
            assign data_11[n746 + d746*16 + c26*28*16] = data_11_array[c26][d746][n746];
        end
    endgenerate
    generate 
        localparam integer d747 = 19;
        for (n747 = 0; n747 < 16; n747 = n747 + 1) 
        begin: outbit747
            assign data_11[n747 + d747*16 + c26*28*16] = data_11_array[c26][d747][n747];
        end
    endgenerate
    generate 
        localparam integer d748 = 20;
        for (n748 = 0; n748 < 16; n748 = n748 + 1) 
        begin: outbit748
            assign data_11[n748 + d748*16 + c26*28*16] = data_11_array[c26][d748][n748];
        end
    endgenerate
    generate 
        localparam integer d749 = 21;
        for (n749 = 0; n749 < 16; n749 = n749 + 1) 
        begin: outbit749
            assign data_11[n749 + d749*16 + c26*28*16] = data_11_array[c26][d749][n749];
        end
    endgenerate
    generate 
        localparam integer d750 = 22;
        for (n750 = 0; n750 < 16; n750 = n750 + 1) 
        begin: outbit750
            assign data_11[n750 + d750*16 + c26*28*16] = data_11_array[c26][d750][n750];
        end
    endgenerate
    generate 
        localparam integer d751 = 23;
        for (n751 = 0; n751 < 16; n751 = n751 + 1) 
        begin: outbit751
            assign data_11[n751 + d751*16 + c26*28*16] = data_11_array[c26][d751][n751];
        end
    endgenerate
    generate 
        localparam integer d752 = 24;
        for (n752 = 0; n752 < 16; n752 = n752 + 1) 
        begin: outbit752
            assign data_11[n752 + d752*16 + c26*28*16] = data_11_array[c26][d752][n752];
        end
    endgenerate
    generate 
        localparam integer d753 = 25;
        for (n753 = 0; n753 < 16; n753 = n753 + 1) 
        begin: outbit753
            assign data_11[n753 + d753*16 + c26*28*16] = data_11_array[c26][d753][n753];
        end
    endgenerate
    generate 
        localparam integer d754 = 26;
        for (n754 = 0; n754 < 16; n754 = n754 + 1) 
        begin: outbit754
            assign data_11[n754 + d754*16 + c26*28*16] = data_11_array[c26][d754][n754];
        end
    endgenerate
    generate 
        localparam integer d755 = 27;
        for (n755 = 0; n755 < 16; n755 = n755 + 1) 
        begin: outbit755
            assign data_11[n755 + d755*16 + c26*28*16] = data_11_array[c26][d755][n755];
        end
    endgenerate
    localparam integer c27 = 27;
    generate 
        localparam integer d756 = 0;
        for (n756 = 0; n756 < 16; n756 = n756 + 1) 
        begin: outbit756
            assign data_11[n756 + d756*16 + c27*28*16] = data_11_array[c27][d756][n756];
        end
    endgenerate
    generate 
        localparam integer d757 = 1;
        for (n757 = 0; n757 < 16; n757 = n757 + 1) 
        begin: outbit757
            assign data_11[n757 + d757*16 + c27*28*16] = data_11_array[c27][d757][n757];
        end
    endgenerate
    generate 
        localparam integer d758 = 2;
        for (n758 = 0; n758 < 16; n758 = n758 + 1) 
        begin: outbit758
            assign data_11[n758 + d758*16 + c27*28*16] = data_11_array[c27][d758][n758];
        end
    endgenerate
    generate 
        localparam integer d759 = 3;
        for (n759 = 0; n759 < 16; n759 = n759 + 1) 
        begin: outbit759
            assign data_11[n759 + d759*16 + c27*28*16] = data_11_array[c27][d759][n759];
        end
    endgenerate
    generate 
        localparam integer d760 = 4;
        for (n760 = 0; n760 < 16; n760 = n760 + 1) 
        begin: outbit760
            assign data_11[n760 + d760*16 + c27*28*16] = data_11_array[c27][d760][n760];
        end
    endgenerate
    generate 
        localparam integer d761 = 5;
        for (n761 = 0; n761 < 16; n761 = n761 + 1) 
        begin: outbit761
            assign data_11[n761 + d761*16 + c27*28*16] = data_11_array[c27][d761][n761];
        end
    endgenerate
    generate 
        localparam integer d762 = 6;
        for (n762 = 0; n762 < 16; n762 = n762 + 1) 
        begin: outbit762
            assign data_11[n762 + d762*16 + c27*28*16] = data_11_array[c27][d762][n762];
        end
    endgenerate
    generate 
        localparam integer d763 = 7;
        for (n763 = 0; n763 < 16; n763 = n763 + 1) 
        begin: outbit763
            assign data_11[n763 + d763*16 + c27*28*16] = data_11_array[c27][d763][n763];
        end
    endgenerate
    generate 
        localparam integer d764 = 8;
        for (n764 = 0; n764 < 16; n764 = n764 + 1) 
        begin: outbit764
            assign data_11[n764 + d764*16 + c27*28*16] = data_11_array[c27][d764][n764];
        end
    endgenerate
    generate 
        localparam integer d765 = 9;
        for (n765 = 0; n765 < 16; n765 = n765 + 1) 
        begin: outbit765
            assign data_11[n765 + d765*16 + c27*28*16] = data_11_array[c27][d765][n765];
        end
    endgenerate
    generate 
        localparam integer d766 = 10;
        for (n766 = 0; n766 < 16; n766 = n766 + 1) 
        begin: outbit766
            assign data_11[n766 + d766*16 + c27*28*16] = data_11_array[c27][d766][n766];
        end
    endgenerate
    generate 
        localparam integer d767 = 11;
        for (n767 = 0; n767 < 16; n767 = n767 + 1) 
        begin: outbit767
            assign data_11[n767 + d767*16 + c27*28*16] = data_11_array[c27][d767][n767];
        end
    endgenerate
    generate 
        localparam integer d768 = 12;
        for (n768 = 0; n768 < 16; n768 = n768 + 1) 
        begin: outbit768
            assign data_11[n768 + d768*16 + c27*28*16] = data_11_array[c27][d768][n768];
        end
    endgenerate
    generate 
        localparam integer d769 = 13;
        for (n769 = 0; n769 < 16; n769 = n769 + 1) 
        begin: outbit769
            assign data_11[n769 + d769*16 + c27*28*16] = data_11_array[c27][d769][n769];
        end
    endgenerate
    generate 
        localparam integer d770 = 14;
        for (n770 = 0; n770 < 16; n770 = n770 + 1) 
        begin: outbit770
            assign data_11[n770 + d770*16 + c27*28*16] = data_11_array[c27][d770][n770];
        end
    endgenerate
    generate 
        localparam integer d771 = 15;
        for (n771 = 0; n771 < 16; n771 = n771 + 1) 
        begin: outbit771
            assign data_11[n771 + d771*16 + c27*28*16] = data_11_array[c27][d771][n771];
        end
    endgenerate
    generate 
        localparam integer d772 = 16;
        for (n772 = 0; n772 < 16; n772 = n772 + 1) 
        begin: outbit772
            assign data_11[n772 + d772*16 + c27*28*16] = data_11_array[c27][d772][n772];
        end
    endgenerate
    generate 
        localparam integer d773 = 17;
        for (n773 = 0; n773 < 16; n773 = n773 + 1) 
        begin: outbit773
            assign data_11[n773 + d773*16 + c27*28*16] = data_11_array[c27][d773][n773];
        end
    endgenerate
    generate 
        localparam integer d774 = 18;
        for (n774 = 0; n774 < 16; n774 = n774 + 1) 
        begin: outbit774
            assign data_11[n774 + d774*16 + c27*28*16] = data_11_array[c27][d774][n774];
        end
    endgenerate
    generate 
        localparam integer d775 = 19;
        for (n775 = 0; n775 < 16; n775 = n775 + 1) 
        begin: outbit775
            assign data_11[n775 + d775*16 + c27*28*16] = data_11_array[c27][d775][n775];
        end
    endgenerate
    generate 
        localparam integer d776 = 20;
        for (n776 = 0; n776 < 16; n776 = n776 + 1) 
        begin: outbit776
            assign data_11[n776 + d776*16 + c27*28*16] = data_11_array[c27][d776][n776];
        end
    endgenerate
    generate 
        localparam integer d777 = 21;
        for (n777 = 0; n777 < 16; n777 = n777 + 1) 
        begin: outbit777
            assign data_11[n777 + d777*16 + c27*28*16] = data_11_array[c27][d777][n777];
        end
    endgenerate
    generate 
        localparam integer d778 = 22;
        for (n778 = 0; n778 < 16; n778 = n778 + 1) 
        begin: outbit778
            assign data_11[n778 + d778*16 + c27*28*16] = data_11_array[c27][d778][n778];
        end
    endgenerate
    generate 
        localparam integer d779 = 23;
        for (n779 = 0; n779 < 16; n779 = n779 + 1) 
        begin: outbit779
            assign data_11[n779 + d779*16 + c27*28*16] = data_11_array[c27][d779][n779];
        end
    endgenerate
    generate 
        localparam integer d780 = 24;
        for (n780 = 0; n780 < 16; n780 = n780 + 1) 
        begin: outbit780
            assign data_11[n780 + d780*16 + c27*28*16] = data_11_array[c27][d780][n780];
        end
    endgenerate
    generate 
        localparam integer d781 = 25;
        for (n781 = 0; n781 < 16; n781 = n781 + 1) 
        begin: outbit781
            assign data_11[n781 + d781*16 + c27*28*16] = data_11_array[c27][d781][n781];
        end
    endgenerate
    generate 
        localparam integer d782 = 26;
        for (n782 = 0; n782 < 16; n782 = n782 + 1) 
        begin: outbit782
            assign data_11[n782 + d782*16 + c27*28*16] = data_11_array[c27][d782][n782];
        end
    endgenerate
    generate 
        localparam integer d783 = 27;
        for (n783 = 0; n783 < 16; n783 = n783 + 1) 
        begin: outbit783
            assign data_11[n783 + d783*16 + c27*28*16] = data_11_array[c27][d783][n783];
        end
    endgenerate
    
endmodule

////CONVOLUTION LAYER 1 | FEATURE MAP 2
module Conv1_feature2 (
    data,
    feature2Weight_0,
    feature2Weight_1,
    feature2Weight_2,
    feature2Weight_3,
    feature2Weight_4,
    feature2Weight_5,
    feature2Weight_6,
    feature2Weight_7,
    feature2Weight_8,
    feature2Weight_9,
    feature2Weight_10,
    feature2Weight_11,
    feature2Weight_12,
    feature2Weight_13,
    feature2Weight_14,
    feature2Weight_15,
    feature2Weight_16,
    feature2Weight_17,
    feature2Weight_18,
    feature2Weight_19,
    feature2Weight_20,
    feature2Weight_21,
    feature2Weight_22,
    feature2Weight_23,
    feature2Weight_24,
    feature2Bias,
    data_11);

  parameter TEST_DATA = 784*16,
    FP_LENGTH = 16;
  input [TEST_DATA - 1:0] data;
  input [FP_LENGTH - 1:0] feature2Weight_0, feature2Weight_1, feature2Weight_2, feature2Weight_3, feature2Weight_4, feature2Weight_5, feature2Weight_6, feature2Weight_7, feature2Weight_8, feature2Weight_9, feature2Weight_10, feature2Weight_11, feature2Weight_12, feature2Weight_13, feature2Weight_14, feature2Weight_15, feature2Weight_16, feature2Weight_17, feature2Weight_18, feature2Weight_19, feature2Weight_20, feature2Weight_21, feature2Weight_22, feature2Weight_23, feature2Weight_24, feature2Bias;
  output [576*16 - 1:0] data_11;    
  
  wire [FP_LENGTH - 1:0] data_array [0:27][0:27];
  wire [FP_LENGTH - 1:0] data_11_array [0:23][0:23];
  wire [FP_LENGTH - 1:0] multi0 [0:24][0:23], multi1 [0:24][0:23], multi2 [0:24][0:23], multi3 [0:24][0:23], multi4 [0:24][0:23], multi5 [0:24][0:23], multi6 [0:24][0:23], multi7 [0:24][0:23], multi8 [0:24][0:23], multi9 [0:24][0:23], multi10 [0:24][0:23], multi11 [0:24][0:23], multi12 [0:24][0:23], multi13 [0:24][0:23], multi14 [0:24][0:23], multi15 [0:24][0:23], multi16 [0:24][0:23], multi17 [0:24][0:23], multi18 [0:24][0:23], multi19 [0:24][0:23], multi20 [0:24][0:23], multi21 [0:24][0:23], multi22 [0:24][0:23], multi23 [0:24][0:23], multi24 [0:24][0:23];
  wire [FP_LENGTH - 1:0] sum0 [0:23][0:23], sum1 [0:23][0:23], sum2 [0:23][0:23], sum3 [0:23][0:23], sum4 [0:23][0:23], sum5 [0:23][0:23], sum6 [0:23][0:23], sum7 [0:23][0:23], sum8 [0:23][0:23], sum9 [0:23][0:23], sum10 [0:23][0:23], sum11 [0:23][0:23], sum12 [0:23][0:23], sum13 [0:23][0:23], sum14 [0:23][0:23], sum15 [0:23][0:23], sum16 [0:23][0:23], sum17 [0:23][0:23], sum18 [0:23][0:23], sum19 [0:23][0:23], sum20 [0:23][0:23], sum21 [0:23][0:23], sum22 [0:23][0:23], sum23 [0:23][0:23], sum24 [0:23][0:23];
//  integer a, b, c; ///a = ROW, b = COLUMN, c = 16 bit Value
  
//  initial begin
//    for (a = 0; a < 28; a = a + 1) begin
//        for (b = 0; b < 28; b = b + 1) begin
//            for (c = 15; c >= 0; c = c - 1) begin
//                data_array[a][b][c] = data[c + b*16 + a*28*16];
//            end
//        end
//    end
    
//    forever begin
//        for (a = 0; a < 28; a = a + 1) begin
//            for (b = 0; b < 28; b = b + 1) begin
//                for (c = 15; c >= 0; c = c - 1) begin
//                   data_11[c + b*16 + a*28*16] = data_11_array[a][b][c];
//                end
//            end
//        end
//    end
//  end
  
  
  
  genvar i0, i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21, i22, i23, i24, m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15,m16,m17,m18,m19,m20,m21,m22,m23,m24,m25,m26,m27,m28,m29,m30,m31,m32,m33,m34,m35,m36,m37,m38,m39,m40,m41,m42,m43,m44,m45,m46,m47,m48,m49,m50,m51,m52,m53,m54,m55,m56,m57,m58,m59,m60,m61,m62,m63,m64,m65,m66,m67,m68,m69,m70,m71,m72,m73,m74,m75,m76,m77,m78,m79,m80,m81,m82,m83,m84,m85,m86,m87,m88,m89,m90,m91,m92,m93,m94,m95,m96,m97,m98,m99,m100,m101,m102,m103,m104,m105,m106,m107,m108,m109,m110,m111,m112,m113,m114,m115,m116,m117,m118,m119,m120,m121,m122,m123,m124,m125,m126,m127,m128,m129,m130,m131,m132,m133,m134,m135,m136,m137,m138,m139,m140,m141,m142,m143,m144,m145,m146,m147,m148,m149,m150,m151,m152,m153,m154,m155,m156,m157,m158,m159,m160,m161,m162,m163,m164,m165,m166,m167,m168,m169,m170,m171,m172,m173,m174,m175,m176,m177,m178,m179,m180,m181,m182,m183,m184,m185,m186,m187,m188,m189,m190,m191,m192,m193,m194,m195,m196,m197,m198,m199,m200,m201,m202,m203,m204,m205,m206,m207,m208,m209,m210,m211,m212,m213,m214,m215,m216,m217,m218,m219,m220,m221,m222,m223,m224,m225,m226,m227,m228,m229,m230,m231,m232,m233,m234,m235,m236,m237,m238,m239,m240,m241,m242,m243,m244,m245,m246,m247,m248,m249,m250,m251,m252,m253,m254,m255,m256,m257,m258,m259,m260,m261,m262,m263,m264,m265,m266,m267,m268,m269,m270,m271,m272,m273,m274,m275,m276,m277,m278,m279,m280,m281,m282,m283,m284,m285,m286,m287,m288,m289,m290,m291,m292,m293,m294,m295,m296,m297,m298,m299,m300,m301,m302,m303,m304,m305,m306,m307,m308,m309,m310,m311,m312,m313,m314,m315,m316,m317,m318,m319,m320,m321,m322,m323,m324,m325,m326,m327,m328,m329,m330,m331,m332,m333,m334,m335,m336,m337,m338,m339,m340,m341,m342,m343,m344,m345,m346,m347,m348,m349,m350,m351,m352,m353,m354,m355,m356,m357,m358,m359,m360,m361,m362,m363,m364,m365,m366,m367,m368,m369,m370,m371,m372,m373,m374,m375,m376,m377,m378,m379,m380,m381,m382,m383,m384,m385,m386,m387,m388,m389,m390,m391,m392,m393,m394,m395,m396,m397,m398,m399,m400,m401,m402,m403,m404,m405,m406,m407,m408,m409,m410,m411,m412,m413,m414,m415,m416,m417,m418,m419,m420,m421,m422,m423,m424,m425,m426,m427,m428,m429,m430,m431,m432,m433,m434,m435,m436,m437,m438,m439,m440,m441,m442,m443,m444,m445,m446,m447,m448,m449,m450,m451,m452,m453,m454,m455,m456,m457,m458,m459,m460,m461,m462,m463,m464,m465,m466,m467,m468,m469,m470,m471,m472,m473,m474,m475,m476,m477,m478,m479,m480,m481,m482,m483,m484,m485,m486,m487,m488,m489,m490,m491,m492,m493,m494,m495,m496,m497,m498,m499,m500,m501,m502,m503,m504,m505,m506,m507,m508,m509,m510,m511,m512,m513,m514,m515,m516,m517,m518,m519,m520,m521,m522,m523,m524,m525,m526,m527,m528,m529,m530,m531,m532,m533,m534,m535,m536,m537,m538,m539,m540,m541,m542,m543,m544,m545,m546,m547,m548,m549,m550,m551,m552,m553,m554,m555,m556,m557,m558,m559,m560,m561,m562,m563,m564,m565,m566,m567,m568,m569,m570,m571,m572,m573,m574,m575,m576,m577,m578,m579,m580,m581,m582,m583,m584,m585,m586,m587,m588,m589,m590,m591,m592,m593,m594,m595,m596,m597,m598,m599,m600,m601,m602,m603,m604,m605,m606,m607,m608,m609,m610,m611,m612,m613,m614,m615,m616,m617,m618,m619,m620,m621,m622,m623,m624,m625,m626,m627,m628,m629,m630,m631,m632,m633,m634,m635,m636,m637,m638,m639,m640,m641,m642,m643,m644,m645,m646,m647,m648,m649,m650,m651,m652,m653,m654,m655,m656,m657,m658,m659,m660,m661,m662,m663,m664,m665,m666,m667,m668,m669,m670,m671,m672,m673,m674,m675,m676,m677,m678,m679,m680,m681,m682,m683,m684,m685,m686,m687,m688,m689,m690,m691,m692,m693,m694,m695,m696,m697,m698,m699,m700,m701,m702,m703,m704,m705,m706,m707,m708,m709,m710,m711,m712,m713,m714,m715,m716,m717,m718,m719,m720,m721,m722,m723,m724,m725,m726,m727,m728,m729,m730,m731,m732,m733,m734,m735,m736,m737,m738,m739,m740,m741,m742,m743,m744,m745,m746,m747,m748,m749,m750,m751,m752,m753,m754,m755,m756,m757,m758,m759,m760,m761,m762,m763,m764,m765,m766,m767,m768,m769,m770,m771,m772,m773,m774,m775,m776,m777,m778,m779,m780,m781,m782,m783,n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n50,n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80,n81,n82,n83,n84,n85,n86,n87,n88,n89,n90,n91,n92,n93,n94,n95,n96,n97,n98,n99,n100,n101,n102,n103,n104,n105,n106,n107,n108,n109,n110,n111,n112,n113,n114,n115,n116,n117,n118,n119,n120,n121,n122,n123,n124,n125,n126,n127,n128,n129,n130,n131,n132,n133,n134,n135,n136,n137,n138,n139,n140,n141,n142,n143,n144,n145,n146,n147,n148,n149,n150,n151,n152,n153,n154,n155,n156,n157,n158,n159,n160,n161,n162,n163,n164,n165,n166,n167,n168,n169,n170,n171,n172,n173,n174,n175,n176,n177,n178,n179,n180,n181,n182,n183,n184,n185,n186,n187,n188,n189,n190,n191,n192,n193,n194,n195,n196,n197,n198,n199,n200,n201,n202,n203,n204,n205,n206,n207,n208,n209,n210,n211,n212,n213,n214,n215,n216,n217,n218,n219,n220,n221,n222,n223,n224,n225,n226,n227,n228,n229,n230,n231,n232,n233,n234,n235,n236,n237,n238,n239,n240,n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,n251,n252,n253,n254,n255,n256,n257,n258,n259,n260,n261,n262,n263,n264,n265,n266,n267,n268,n269,n270,n271,n272,n273,n274,n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,n330,n331,n332,n333,n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,n345,n346,n347,n348,n349,n350,n351,n352,n353,n354,n355,n356,n357,n358,n359,n360,n361,n362,n363,n364,n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,n385,n386,n387,n388,n389,n390,n391,n392,n393,n394,n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,n415,n416,n417,n418,n419,n420,n421,n422,n423,n424,n425,n426,n427,n428,n429,n430,n431,n432,n433,n434,n435,n436,n437,n438,n439,n440,n441,n442,n443,n444,n445,n446,n447,n448,n449,n450,n451,n452,n453,n454,n455,n456,n457,n458,n459,n460,n461,n462,n463,n464,n465,n466,n467,n468,n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,n479,n480,n481,n482,n483,n484,n485,n486,n487,n488,n489,n490,n491,n492,n493,n494,n495,n496,n497,n498,n499,n500,n501,n502,n503,n504,n505,n506,n507,n508,n509,n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,n559,n560,n561,n562,n563,n564,n565,n566,n567,n568,n569,n570,n571,n572,n573,n574,n575,n576,n577,n578,n579,n580,n581,n582,n583,n584,n585,n586,n587,n588,n589,n590,n591,n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,n612,n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,n623,n624,n625,n626,n627,n628,n629,n630,n631,n632,n633,n634,n635,n636,n637,n638,n639,n640,n641,n642,n643,n644,n645,n646,n647,n648,n649,n650,n651,n652,n653,n654,n655,n656,n657,n658,n659,n660,n661,n662,n663,n664,n665,n666,n667,n668,n669,n670,n671,n672,n673,n674,n675,n676,n677,n678,n679,n680,n681,n682,n683,n684,n685,n686,n687,n688,n689,n690,n691,n692,n693,n694,n695,n696,n697,n698,n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,n709,n710,n711,n712,n713,n714,n715,n716,n717,n718,n719,n720,n721,n722,n723,n724,n725,n726,n727,n728,n729,n730,n731,n732,n733,n734,n735,n736,n737,n738,n739,n740,n741,n742,n743,n744,n745,n746,n747,n748,n749,n750,n751,n752,n753,n754,n755,n756,n757,n758,n759,n760,n761,n762,n763,n764,n765,n766,n767,n768,n769,n770,n771,n772,n773,n774,n775,n776,n777,n778,n779,n780,n781,n782,n783;
  
  localparam integer a0 = 0;
    generate 
        localparam integer b0 = 0;
        for (m0 = 0; m0 < 16; m0 = m0 + 1) 
        begin: inbit0
            assign data_11[m0 + b0*16 + a0*28*16] = data_11_array[a0][b0][m0];
        end
    endgenerate
    generate 
        localparam integer b1 = 1;
        for (m1 = 0; m1 < 16; m1 = m1 + 1) 
        begin: inbit1
            assign data_11[m1 + b1*16 + a0*28*16] = data_11_array[a0][b1][m1];
        end
    endgenerate
    generate 
        localparam integer b2 = 2;
        for (m2 = 0; m2 < 16; m2 = m2 + 1) 
        begin: inbit2
            assign data_11[m2 + b2*16 + a0*28*16] = data_11_array[a0][b2][m2];
        end
    endgenerate
    generate 
        localparam integer b3 = 3;
        for (m3 = 0; m3 < 16; m3 = m3 + 1) 
        begin: inbit3
            assign data_11[m3 + b3*16 + a0*28*16] = data_11_array[a0][b3][m3];
        end
    endgenerate
    generate 
        localparam integer b4 = 4;
        for (m4 = 0; m4 < 16; m4 = m4 + 1) 
        begin: inbit4
            assign data_11[m4 + b4*16 + a0*28*16] = data_11_array[a0][b4][m4];
        end
    endgenerate
    generate 
        localparam integer b5 = 5;
        for (m5 = 0; m5 < 16; m5 = m5 + 1) 
        begin: inbit5
            assign data_11[m5 + b5*16 + a0*28*16] = data_11_array[a0][b5][m5];
        end
    endgenerate
    generate 
        localparam integer b6 = 6;
        for (m6 = 0; m6 < 16; m6 = m6 + 1) 
        begin: inbit6
            assign data_11[m6 + b6*16 + a0*28*16] = data_11_array[a0][b6][m6];
        end
    endgenerate
    generate 
        localparam integer b7 = 7;
        for (m7 = 0; m7 < 16; m7 = m7 + 1) 
        begin: inbit7
            assign data_11[m7 + b7*16 + a0*28*16] = data_11_array[a0][b7][m7];
        end
    endgenerate
    generate 
        localparam integer b8 = 8;
        for (m8 = 0; m8 < 16; m8 = m8 + 1) 
        begin: inbit8
            assign data_11[m8 + b8*16 + a0*28*16] = data_11_array[a0][b8][m8];
        end
    endgenerate
    generate 
        localparam integer b9 = 9;
        for (m9 = 0; m9 < 16; m9 = m9 + 1) 
        begin: inbit9
            assign data_11[m9 + b9*16 + a0*28*16] = data_11_array[a0][b9][m9];
        end
    endgenerate
    generate 
        localparam integer b10 = 10;
        for (m10 = 0; m10 < 16; m10 = m10 + 1) 
        begin: inbit10
            assign data_11[m10 + b10*16 + a0*28*16] = data_11_array[a0][b10][m10];
        end
    endgenerate
    generate 
        localparam integer b11 = 11;
        for (m11 = 0; m11 < 16; m11 = m11 + 1) 
        begin: inbit11
            assign data_11[m11 + b11*16 + a0*28*16] = data_11_array[a0][b11][m11];
        end
    endgenerate
    generate 
        localparam integer b12 = 12;
        for (m12 = 0; m12 < 16; m12 = m12 + 1) 
        begin: inbit12
            assign data_11[m12 + b12*16 + a0*28*16] = data_11_array[a0][b12][m12];
        end
    endgenerate
    generate 
        localparam integer b13 = 13;
        for (m13 = 0; m13 < 16; m13 = m13 + 1) 
        begin: inbit13
            assign data_11[m13 + b13*16 + a0*28*16] = data_11_array[a0][b13][m13];
        end
    endgenerate
    generate 
        localparam integer b14 = 14;
        for (m14 = 0; m14 < 16; m14 = m14 + 1) 
        begin: inbit14
            assign data_11[m14 + b14*16 + a0*28*16] = data_11_array[a0][b14][m14];
        end
    endgenerate
    generate 
        localparam integer b15 = 15;
        for (m15 = 0; m15 < 16; m15 = m15 + 1) 
        begin: inbit15
            assign data_11[m15 + b15*16 + a0*28*16] = data_11_array[a0][b15][m15];
        end
    endgenerate
    generate 
        localparam integer b16 = 16;
        for (m16 = 0; m16 < 16; m16 = m16 + 1) 
        begin: inbit16
            assign data_11[m16 + b16*16 + a0*28*16] = data_11_array[a0][b16][m16];
        end
    endgenerate
    generate 
        localparam integer b17 = 17;
        for (m17 = 0; m17 < 16; m17 = m17 + 1) 
        begin: inbit17
            assign data_11[m17 + b17*16 + a0*28*16] = data_11_array[a0][b17][m17];
        end
    endgenerate
    generate 
        localparam integer b18 = 18;
        for (m18 = 0; m18 < 16; m18 = m18 + 1) 
        begin: inbit18
            assign data_11[m18 + b18*16 + a0*28*16] = data_11_array[a0][b18][m18];
        end
    endgenerate
    generate 
        localparam integer b19 = 19;
        for (m19 = 0; m19 < 16; m19 = m19 + 1) 
        begin: inbit19
            assign data_11[m19 + b19*16 + a0*28*16] = data_11_array[a0][b19][m19];
        end
    endgenerate
    generate 
        localparam integer b20 = 20;
        for (m20 = 0; m20 < 16; m20 = m20 + 1) 
        begin: inbit20
            assign data_11[m20 + b20*16 + a0*28*16] = data_11_array[a0][b20][m20];
        end
    endgenerate
    generate 
        localparam integer b21 = 21;
        for (m21 = 0; m21 < 16; m21 = m21 + 1) 
        begin: inbit21
            assign data_11[m21 + b21*16 + a0*28*16] = data_11_array[a0][b21][m21];
        end
    endgenerate
    generate 
        localparam integer b22 = 22;
        for (m22 = 0; m22 < 16; m22 = m22 + 1) 
        begin: inbit22
            assign data_11[m22 + b22*16 + a0*28*16] = data_11_array[a0][b22][m22];
        end
    endgenerate
    generate 
        localparam integer b23 = 23;
        for (m23 = 0; m23 < 16; m23 = m23 + 1) 
        begin: inbit23
            assign data_11[m23 + b23*16 + a0*28*16] = data_11_array[a0][b23][m23];
        end
    endgenerate
    generate 
        localparam integer b24 = 24;
        for (m24 = 0; m24 < 16; m24 = m24 + 1) 
        begin: inbit24
            assign data_11[m24 + b24*16 + a0*28*16] = data_11_array[a0][b24][m24];
        end
    endgenerate
    generate 
        localparam integer b25 = 25;
        for (m25 = 0; m25 < 16; m25 = m25 + 1) 
        begin: inbit25
            assign data_11[m25 + b25*16 + a0*28*16] = data_11_array[a0][b25][m25];
        end
    endgenerate
    generate 
        localparam integer b26 = 26;
        for (m26 = 0; m26 < 16; m26 = m26 + 1) 
        begin: inbit26
            assign data_11[m26 + b26*16 + a0*28*16] = data_11_array[a0][b26][m26];
        end
    endgenerate
    generate 
        localparam integer b27 = 27;
        for (m27 = 0; m27 < 16; m27 = m27 + 1) 
        begin: inbit27
            assign data_11[m27 + b27*16 + a0*28*16] = data_11_array[a0][b27][m27];
        end
    endgenerate
    localparam integer a1 = 1;
    generate 
        localparam integer b28 = 0;
        for (m28 = 0; m28 < 16; m28 = m28 + 1) 
        begin: inbit28
            assign data_11[m28 + b28*16 + a1*28*16] = data_11_array[a1][b28][m28];
        end
    endgenerate
    generate 
        localparam integer b29 = 1;
        for (m29 = 0; m29 < 16; m29 = m29 + 1) 
        begin: inbit29
            assign data_11[m29 + b29*16 + a1*28*16] = data_11_array[a1][b29][m29];
        end
    endgenerate
    generate 
        localparam integer b30 = 2;
        for (m30 = 0; m30 < 16; m30 = m30 + 1) 
        begin: inbit30
            assign data_11[m30 + b30*16 + a1*28*16] = data_11_array[a1][b30][m30];
        end
    endgenerate
    generate 
        localparam integer b31 = 3;
        for (m31 = 0; m31 < 16; m31 = m31 + 1) 
        begin: inbit31
            assign data_11[m31 + b31*16 + a1*28*16] = data_11_array[a1][b31][m31];
        end
    endgenerate
    generate 
        localparam integer b32 = 4;
        for (m32 = 0; m32 < 16; m32 = m32 + 1) 
        begin: inbit32
            assign data_11[m32 + b32*16 + a1*28*16] = data_11_array[a1][b32][m32];
        end
    endgenerate
    generate 
        localparam integer b33 = 5;
        for (m33 = 0; m33 < 16; m33 = m33 + 1) 
        begin: inbit33
            assign data_11[m33 + b33*16 + a1*28*16] = data_11_array[a1][b33][m33];
        end
    endgenerate
    generate 
        localparam integer b34 = 6;
        for (m34 = 0; m34 < 16; m34 = m34 + 1) 
        begin: inbit34
            assign data_11[m34 + b34*16 + a1*28*16] = data_11_array[a1][b34][m34];
        end
    endgenerate
    generate 
        localparam integer b35 = 7;
        for (m35 = 0; m35 < 16; m35 = m35 + 1) 
        begin: inbit35
            assign data_11[m35 + b35*16 + a1*28*16] = data_11_array[a1][b35][m35];
        end
    endgenerate
    generate 
        localparam integer b36 = 8;
        for (m36 = 0; m36 < 16; m36 = m36 + 1) 
        begin: inbit36
            assign data_11[m36 + b36*16 + a1*28*16] = data_11_array[a1][b36][m36];
        end
    endgenerate
    generate 
        localparam integer b37 = 9;
        for (m37 = 0; m37 < 16; m37 = m37 + 1) 
        begin: inbit37
            assign data_11[m37 + b37*16 + a1*28*16] = data_11_array[a1][b37][m37];
        end
    endgenerate
    generate 
        localparam integer b38 = 10;
        for (m38 = 0; m38 < 16; m38 = m38 + 1) 
        begin: inbit38
            assign data_11[m38 + b38*16 + a1*28*16] = data_11_array[a1][b38][m38];
        end
    endgenerate
    generate 
        localparam integer b39 = 11;
        for (m39 = 0; m39 < 16; m39 = m39 + 1) 
        begin: inbit39
            assign data_11[m39 + b39*16 + a1*28*16] = data_11_array[a1][b39][m39];
        end
    endgenerate
    generate 
        localparam integer b40 = 12;
        for (m40 = 0; m40 < 16; m40 = m40 + 1) 
        begin: inbit40
            assign data_11[m40 + b40*16 + a1*28*16] = data_11_array[a1][b40][m40];
        end
    endgenerate
    generate 
        localparam integer b41 = 13;
        for (m41 = 0; m41 < 16; m41 = m41 + 1) 
        begin: inbit41
            assign data_11[m41 + b41*16 + a1*28*16] = data_11_array[a1][b41][m41];
        end
    endgenerate
    generate 
        localparam integer b42 = 14;
        for (m42 = 0; m42 < 16; m42 = m42 + 1) 
        begin: inbit42
            assign data_11[m42 + b42*16 + a1*28*16] = data_11_array[a1][b42][m42];
        end
    endgenerate
    generate 
        localparam integer b43 = 15;
        for (m43 = 0; m43 < 16; m43 = m43 + 1) 
        begin: inbit43
            assign data_11[m43 + b43*16 + a1*28*16] = data_11_array[a1][b43][m43];
        end
    endgenerate
    generate 
        localparam integer b44 = 16;
        for (m44 = 0; m44 < 16; m44 = m44 + 1) 
        begin: inbit44
            assign data_11[m44 + b44*16 + a1*28*16] = data_11_array[a1][b44][m44];
        end
    endgenerate
    generate 
        localparam integer b45 = 17;
        for (m45 = 0; m45 < 16; m45 = m45 + 1) 
        begin: inbit45
            assign data_11[m45 + b45*16 + a1*28*16] = data_11_array[a1][b45][m45];
        end
    endgenerate
    generate 
        localparam integer b46 = 18;
        for (m46 = 0; m46 < 16; m46 = m46 + 1) 
        begin: inbit46
            assign data_11[m46 + b46*16 + a1*28*16] = data_11_array[a1][b46][m46];
        end
    endgenerate
    generate 
        localparam integer b47 = 19;
        for (m47 = 0; m47 < 16; m47 = m47 + 1) 
        begin: inbit47
            assign data_11[m47 + b47*16 + a1*28*16] = data_11_array[a1][b47][m47];
        end
    endgenerate
    generate 
        localparam integer b48 = 20;
        for (m48 = 0; m48 < 16; m48 = m48 + 1) 
        begin: inbit48
            assign data_11[m48 + b48*16 + a1*28*16] = data_11_array[a1][b48][m48];
        end
    endgenerate
    generate 
        localparam integer b49 = 21;
        for (m49 = 0; m49 < 16; m49 = m49 + 1) 
        begin: inbit49
            assign data_11[m49 + b49*16 + a1*28*16] = data_11_array[a1][b49][m49];
        end
    endgenerate
    generate 
        localparam integer b50 = 22;
        for (m50 = 0; m50 < 16; m50 = m50 + 1) 
        begin: inbit50
            assign data_11[m50 + b50*16 + a1*28*16] = data_11_array[a1][b50][m50];
        end
    endgenerate
    generate 
        localparam integer b51 = 23;
        for (m51 = 0; m51 < 16; m51 = m51 + 1) 
        begin: inbit51
            assign data_11[m51 + b51*16 + a1*28*16] = data_11_array[a1][b51][m51];
        end
    endgenerate
    generate 
        localparam integer b52 = 24;
        for (m52 = 0; m52 < 16; m52 = m52 + 1) 
        begin: inbit52
            assign data_11[m52 + b52*16 + a1*28*16] = data_11_array[a1][b52][m52];
        end
    endgenerate
    generate 
        localparam integer b53 = 25;
        for (m53 = 0; m53 < 16; m53 = m53 + 1) 
        begin: inbit53
            assign data_11[m53 + b53*16 + a1*28*16] = data_11_array[a1][b53][m53];
        end
    endgenerate
    generate 
        localparam integer b54 = 26;
        for (m54 = 0; m54 < 16; m54 = m54 + 1) 
        begin: inbit54
            assign data_11[m54 + b54*16 + a1*28*16] = data_11_array[a1][b54][m54];
        end
    endgenerate
    generate 
        localparam integer b55 = 27;
        for (m55 = 0; m55 < 16; m55 = m55 + 1) 
        begin: inbit55
            assign data_11[m55 + b55*16 + a1*28*16] = data_11_array[a1][b55][m55];
        end
    endgenerate
    localparam integer a2 = 2;
    generate 
        localparam integer b56 = 0;
        for (m56 = 0; m56 < 16; m56 = m56 + 1) 
        begin: inbit56
            assign data_11[m56 + b56*16 + a2*28*16] = data_11_array[a2][b56][m56];
        end
    endgenerate
    generate 
        localparam integer b57 = 1;
        for (m57 = 0; m57 < 16; m57 = m57 + 1) 
        begin: inbit57
            assign data_11[m57 + b57*16 + a2*28*16] = data_11_array[a2][b57][m57];
        end
    endgenerate
    generate 
        localparam integer b58 = 2;
        for (m58 = 0; m58 < 16; m58 = m58 + 1) 
        begin: inbit58
            assign data_11[m58 + b58*16 + a2*28*16] = data_11_array[a2][b58][m58];
        end
    endgenerate
    generate 
        localparam integer b59 = 3;
        for (m59 = 0; m59 < 16; m59 = m59 + 1) 
        begin: inbit59
            assign data_11[m59 + b59*16 + a2*28*16] = data_11_array[a2][b59][m59];
        end
    endgenerate
    generate 
        localparam integer b60 = 4;
        for (m60 = 0; m60 < 16; m60 = m60 + 1) 
        begin: inbit60
            assign data_11[m60 + b60*16 + a2*28*16] = data_11_array[a2][b60][m60];
        end
    endgenerate
    generate 
        localparam integer b61 = 5;
        for (m61 = 0; m61 < 16; m61 = m61 + 1) 
        begin: inbit61
            assign data_11[m61 + b61*16 + a2*28*16] = data_11_array[a2][b61][m61];
        end
    endgenerate
    generate 
        localparam integer b62 = 6;
        for (m62 = 0; m62 < 16; m62 = m62 + 1) 
        begin: inbit62
            assign data_11[m62 + b62*16 + a2*28*16] = data_11_array[a2][b62][m62];
        end
    endgenerate
    generate 
        localparam integer b63 = 7;
        for (m63 = 0; m63 < 16; m63 = m63 + 1) 
        begin: inbit63
            assign data_11[m63 + b63*16 + a2*28*16] = data_11_array[a2][b63][m63];
        end
    endgenerate
    generate 
        localparam integer b64 = 8;
        for (m64 = 0; m64 < 16; m64 = m64 + 1) 
        begin: inbit64
            assign data_11[m64 + b64*16 + a2*28*16] = data_11_array[a2][b64][m64];
        end
    endgenerate
    generate 
        localparam integer b65 = 9;
        for (m65 = 0; m65 < 16; m65 = m65 + 1) 
        begin: inbit65
            assign data_11[m65 + b65*16 + a2*28*16] = data_11_array[a2][b65][m65];
        end
    endgenerate
    generate 
        localparam integer b66 = 10;
        for (m66 = 0; m66 < 16; m66 = m66 + 1) 
        begin: inbit66
            assign data_11[m66 + b66*16 + a2*28*16] = data_11_array[a2][b66][m66];
        end
    endgenerate
    generate 
        localparam integer b67 = 11;
        for (m67 = 0; m67 < 16; m67 = m67 + 1) 
        begin: inbit67
            assign data_11[m67 + b67*16 + a2*28*16] = data_11_array[a2][b67][m67];
        end
    endgenerate
    generate 
        localparam integer b68 = 12;
        for (m68 = 0; m68 < 16; m68 = m68 + 1) 
        begin: inbit68
            assign data_11[m68 + b68*16 + a2*28*16] = data_11_array[a2][b68][m68];
        end
    endgenerate
    generate 
        localparam integer b69 = 13;
        for (m69 = 0; m69 < 16; m69 = m69 + 1) 
        begin: inbit69
            assign data_11[m69 + b69*16 + a2*28*16] = data_11_array[a2][b69][m69];
        end
    endgenerate
    generate 
        localparam integer b70 = 14;
        for (m70 = 0; m70 < 16; m70 = m70 + 1) 
        begin: inbit70
            assign data_11[m70 + b70*16 + a2*28*16] = data_11_array[a2][b70][m70];
        end
    endgenerate
    generate 
        localparam integer b71 = 15;
        for (m71 = 0; m71 < 16; m71 = m71 + 1) 
        begin: inbit71
            assign data_11[m71 + b71*16 + a2*28*16] = data_11_array[a2][b71][m71];
        end
    endgenerate
    generate 
        localparam integer b72 = 16;
        for (m72 = 0; m72 < 16; m72 = m72 + 1) 
        begin: inbit72
            assign data_11[m72 + b72*16 + a2*28*16] = data_11_array[a2][b72][m72];
        end
    endgenerate
    generate 
        localparam integer b73 = 17;
        for (m73 = 0; m73 < 16; m73 = m73 + 1) 
        begin: inbit73
            assign data_11[m73 + b73*16 + a2*28*16] = data_11_array[a2][b73][m73];
        end
    endgenerate
    generate 
        localparam integer b74 = 18;
        for (m74 = 0; m74 < 16; m74 = m74 + 1) 
        begin: inbit74
            assign data_11[m74 + b74*16 + a2*28*16] = data_11_array[a2][b74][m74];
        end
    endgenerate
    generate 
        localparam integer b75 = 19;
        for (m75 = 0; m75 < 16; m75 = m75 + 1) 
        begin: inbit75
            assign data_11[m75 + b75*16 + a2*28*16] = data_11_array[a2][b75][m75];
        end
    endgenerate
    generate 
        localparam integer b76 = 20;
        for (m76 = 0; m76 < 16; m76 = m76 + 1) 
        begin: inbit76
            assign data_11[m76 + b76*16 + a2*28*16] = data_11_array[a2][b76][m76];
        end
    endgenerate
    generate 
        localparam integer b77 = 21;
        for (m77 = 0; m77 < 16; m77 = m77 + 1) 
        begin: inbit77
            assign data_11[m77 + b77*16 + a2*28*16] = data_11_array[a2][b77][m77];
        end
    endgenerate
    generate 
        localparam integer b78 = 22;
        for (m78 = 0; m78 < 16; m78 = m78 + 1) 
        begin: inbit78
            assign data_11[m78 + b78*16 + a2*28*16] = data_11_array[a2][b78][m78];
        end
    endgenerate
    generate 
        localparam integer b79 = 23;
        for (m79 = 0; m79 < 16; m79 = m79 + 1) 
        begin: inbit79
            assign data_11[m79 + b79*16 + a2*28*16] = data_11_array[a2][b79][m79];
        end
    endgenerate
    generate 
        localparam integer b80 = 24;
        for (m80 = 0; m80 < 16; m80 = m80 + 1) 
        begin: inbit80
            assign data_11[m80 + b80*16 + a2*28*16] = data_11_array[a2][b80][m80];
        end
    endgenerate
    generate 
        localparam integer b81 = 25;
        for (m81 = 0; m81 < 16; m81 = m81 + 1) 
        begin: inbit81
            assign data_11[m81 + b81*16 + a2*28*16] = data_11_array[a2][b81][m81];
        end
    endgenerate
    generate 
        localparam integer b82 = 26;
        for (m82 = 0; m82 < 16; m82 = m82 + 1) 
        begin: inbit82
            assign data_11[m82 + b82*16 + a2*28*16] = data_11_array[a2][b82][m82];
        end
    endgenerate
    generate 
        localparam integer b83 = 27;
        for (m83 = 0; m83 < 16; m83 = m83 + 1) 
        begin: inbit83
            assign data_11[m83 + b83*16 + a2*28*16] = data_11_array[a2][b83][m83];
        end
    endgenerate
    localparam integer a3 = 3;
    generate 
        localparam integer b84 = 0;
        for (m84 = 0; m84 < 16; m84 = m84 + 1) 
        begin: inbit84
            assign data_11[m84 + b84*16 + a3*28*16] = data_11_array[a3][b84][m84];
        end
    endgenerate
    generate 
        localparam integer b85 = 1;
        for (m85 = 0; m85 < 16; m85 = m85 + 1) 
        begin: inbit85
            assign data_11[m85 + b85*16 + a3*28*16] = data_11_array[a3][b85][m85];
        end
    endgenerate
    generate 
        localparam integer b86 = 2;
        for (m86 = 0; m86 < 16; m86 = m86 + 1) 
        begin: inbit86
            assign data_11[m86 + b86*16 + a3*28*16] = data_11_array[a3][b86][m86];
        end
    endgenerate
    generate 
        localparam integer b87 = 3;
        for (m87 = 0; m87 < 16; m87 = m87 + 1) 
        begin: inbit87
            assign data_11[m87 + b87*16 + a3*28*16] = data_11_array[a3][b87][m87];
        end
    endgenerate
    generate 
        localparam integer b88 = 4;
        for (m88 = 0; m88 < 16; m88 = m88 + 1) 
        begin: inbit88
            assign data_11[m88 + b88*16 + a3*28*16] = data_11_array[a3][b88][m88];
        end
    endgenerate
    generate 
        localparam integer b89 = 5;
        for (m89 = 0; m89 < 16; m89 = m89 + 1) 
        begin: inbit89
            assign data_11[m89 + b89*16 + a3*28*16] = data_11_array[a3][b89][m89];
        end
    endgenerate
    generate 
        localparam integer b90 = 6;
        for (m90 = 0; m90 < 16; m90 = m90 + 1) 
        begin: inbit90
            assign data_11[m90 + b90*16 + a3*28*16] = data_11_array[a3][b90][m90];
        end
    endgenerate
    generate 
        localparam integer b91 = 7;
        for (m91 = 0; m91 < 16; m91 = m91 + 1) 
        begin: inbit91
            assign data_11[m91 + b91*16 + a3*28*16] = data_11_array[a3][b91][m91];
        end
    endgenerate
    generate 
        localparam integer b92 = 8;
        for (m92 = 0; m92 < 16; m92 = m92 + 1) 
        begin: inbit92
            assign data_11[m92 + b92*16 + a3*28*16] = data_11_array[a3][b92][m92];
        end
    endgenerate
    generate 
        localparam integer b93 = 9;
        for (m93 = 0; m93 < 16; m93 = m93 + 1) 
        begin: inbit93
            assign data_11[m93 + b93*16 + a3*28*16] = data_11_array[a3][b93][m93];
        end
    endgenerate
    generate 
        localparam integer b94 = 10;
        for (m94 = 0; m94 < 16; m94 = m94 + 1) 
        begin: inbit94
            assign data_11[m94 + b94*16 + a3*28*16] = data_11_array[a3][b94][m94];
        end
    endgenerate
    generate 
        localparam integer b95 = 11;
        for (m95 = 0; m95 < 16; m95 = m95 + 1) 
        begin: inbit95
            assign data_11[m95 + b95*16 + a3*28*16] = data_11_array[a3][b95][m95];
        end
    endgenerate
    generate 
        localparam integer b96 = 12;
        for (m96 = 0; m96 < 16; m96 = m96 + 1) 
        begin: inbit96
            assign data_11[m96 + b96*16 + a3*28*16] = data_11_array[a3][b96][m96];
        end
    endgenerate
    generate 
        localparam integer b97 = 13;
        for (m97 = 0; m97 < 16; m97 = m97 + 1) 
        begin: inbit97
            assign data_11[m97 + b97*16 + a3*28*16] = data_11_array[a3][b97][m97];
        end
    endgenerate
    generate 
        localparam integer b98 = 14;
        for (m98 = 0; m98 < 16; m98 = m98 + 1) 
        begin: inbit98
            assign data_11[m98 + b98*16 + a3*28*16] = data_11_array[a3][b98][m98];
        end
    endgenerate
    generate 
        localparam integer b99 = 15;
        for (m99 = 0; m99 < 16; m99 = m99 + 1) 
        begin: inbit99
            assign data_11[m99 + b99*16 + a3*28*16] = data_11_array[a3][b99][m99];
        end
    endgenerate
    generate 
        localparam integer b100 = 16;
        for (m100 = 0; m100 < 16; m100 = m100 + 1) 
        begin: inbit100
            assign data_11[m100 + b100*16 + a3*28*16] = data_11_array[a3][b100][m100];
        end
    endgenerate
    generate 
        localparam integer b101 = 17;
        for (m101 = 0; m101 < 16; m101 = m101 + 1) 
        begin: inbit101
            assign data_11[m101 + b101*16 + a3*28*16] = data_11_array[a3][b101][m101];
        end
    endgenerate
    generate 
        localparam integer b102 = 18;
        for (m102 = 0; m102 < 16; m102 = m102 + 1) 
        begin: inbit102
            assign data_11[m102 + b102*16 + a3*28*16] = data_11_array[a3][b102][m102];
        end
    endgenerate
    generate 
        localparam integer b103 = 19;
        for (m103 = 0; m103 < 16; m103 = m103 + 1) 
        begin: inbit103
            assign data_11[m103 + b103*16 + a3*28*16] = data_11_array[a3][b103][m103];
        end
    endgenerate
    generate 
        localparam integer b104 = 20;
        for (m104 = 0; m104 < 16; m104 = m104 + 1) 
        begin: inbit104
            assign data_11[m104 + b104*16 + a3*28*16] = data_11_array[a3][b104][m104];
        end
    endgenerate
    generate 
        localparam integer b105 = 21;
        for (m105 = 0; m105 < 16; m105 = m105 + 1) 
        begin: inbit105
            assign data_11[m105 + b105*16 + a3*28*16] = data_11_array[a3][b105][m105];
        end
    endgenerate
    generate 
        localparam integer b106 = 22;
        for (m106 = 0; m106 < 16; m106 = m106 + 1) 
        begin: inbit106
            assign data_11[m106 + b106*16 + a3*28*16] = data_11_array[a3][b106][m106];
        end
    endgenerate
    generate 
        localparam integer b107 = 23;
        for (m107 = 0; m107 < 16; m107 = m107 + 1) 
        begin: inbit107
            assign data_11[m107 + b107*16 + a3*28*16] = data_11_array[a3][b107][m107];
        end
    endgenerate
    generate 
        localparam integer b108 = 24;
        for (m108 = 0; m108 < 16; m108 = m108 + 1) 
        begin: inbit108
            assign data_11[m108 + b108*16 + a3*28*16] = data_11_array[a3][b108][m108];
        end
    endgenerate
    generate 
        localparam integer b109 = 25;
        for (m109 = 0; m109 < 16; m109 = m109 + 1) 
        begin: inbit109
            assign data_11[m109 + b109*16 + a3*28*16] = data_11_array[a3][b109][m109];
        end
    endgenerate
    generate 
        localparam integer b110 = 26;
        for (m110 = 0; m110 < 16; m110 = m110 + 1) 
        begin: inbit110
            assign data_11[m110 + b110*16 + a3*28*16] = data_11_array[a3][b110][m110];
        end
    endgenerate
    generate 
        localparam integer b111 = 27;
        for (m111 = 0; m111 < 16; m111 = m111 + 1) 
        begin: inbit111
            assign data_11[m111 + b111*16 + a3*28*16] = data_11_array[a3][b111][m111];
        end
    endgenerate
    localparam integer a4 = 4;
    generate 
        localparam integer b112 = 0;
        for (m112 = 0; m112 < 16; m112 = m112 + 1) 
        begin: inbit112
            assign data_11[m112 + b112*16 + a4*28*16] = data_11_array[a4][b112][m112];
        end
    endgenerate
    generate 
        localparam integer b113 = 1;
        for (m113 = 0; m113 < 16; m113 = m113 + 1) 
        begin: inbit113
            assign data_11[m113 + b113*16 + a4*28*16] = data_11_array[a4][b113][m113];
        end
    endgenerate
    generate 
        localparam integer b114 = 2;
        for (m114 = 0; m114 < 16; m114 = m114 + 1) 
        begin: inbit114
            assign data_11[m114 + b114*16 + a4*28*16] = data_11_array[a4][b114][m114];
        end
    endgenerate
    generate 
        localparam integer b115 = 3;
        for (m115 = 0; m115 < 16; m115 = m115 + 1) 
        begin: inbit115
            assign data_11[m115 + b115*16 + a4*28*16] = data_11_array[a4][b115][m115];
        end
    endgenerate
    generate 
        localparam integer b116 = 4;
        for (m116 = 0; m116 < 16; m116 = m116 + 1) 
        begin: inbit116
            assign data_11[m116 + b116*16 + a4*28*16] = data_11_array[a4][b116][m116];
        end
    endgenerate
    generate 
        localparam integer b117 = 5;
        for (m117 = 0; m117 < 16; m117 = m117 + 1) 
        begin: inbit117
            assign data_11[m117 + b117*16 + a4*28*16] = data_11_array[a4][b117][m117];
        end
    endgenerate
    generate 
        localparam integer b118 = 6;
        for (m118 = 0; m118 < 16; m118 = m118 + 1) 
        begin: inbit118
            assign data_11[m118 + b118*16 + a4*28*16] = data_11_array[a4][b118][m118];
        end
    endgenerate
    generate 
        localparam integer b119 = 7;
        for (m119 = 0; m119 < 16; m119 = m119 + 1) 
        begin: inbit119
            assign data_11[m119 + b119*16 + a4*28*16] = data_11_array[a4][b119][m119];
        end
    endgenerate
    generate 
        localparam integer b120 = 8;
        for (m120 = 0; m120 < 16; m120 = m120 + 1) 
        begin: inbit120
            assign data_11[m120 + b120*16 + a4*28*16] = data_11_array[a4][b120][m120];
        end
    endgenerate
    generate 
        localparam integer b121 = 9;
        for (m121 = 0; m121 < 16; m121 = m121 + 1) 
        begin: inbit121
            assign data_11[m121 + b121*16 + a4*28*16] = data_11_array[a4][b121][m121];
        end
    endgenerate
    generate 
        localparam integer b122 = 10;
        for (m122 = 0; m122 < 16; m122 = m122 + 1) 
        begin: inbit122
            assign data_11[m122 + b122*16 + a4*28*16] = data_11_array[a4][b122][m122];
        end
    endgenerate
    generate 
        localparam integer b123 = 11;
        for (m123 = 0; m123 < 16; m123 = m123 + 1) 
        begin: inbit123
            assign data_11[m123 + b123*16 + a4*28*16] = data_11_array[a4][b123][m123];
        end
    endgenerate
    generate 
        localparam integer b124 = 12;
        for (m124 = 0; m124 < 16; m124 = m124 + 1) 
        begin: inbit124
            assign data_11[m124 + b124*16 + a4*28*16] = data_11_array[a4][b124][m124];
        end
    endgenerate
    generate 
        localparam integer b125 = 13;
        for (m125 = 0; m125 < 16; m125 = m125 + 1) 
        begin: inbit125
            assign data_11[m125 + b125*16 + a4*28*16] = data_11_array[a4][b125][m125];
        end
    endgenerate
    generate 
        localparam integer b126 = 14;
        for (m126 = 0; m126 < 16; m126 = m126 + 1) 
        begin: inbit126
            assign data_11[m126 + b126*16 + a4*28*16] = data_11_array[a4][b126][m126];
        end
    endgenerate
    generate 
        localparam integer b127 = 15;
        for (m127 = 0; m127 < 16; m127 = m127 + 1) 
        begin: inbit127
            assign data_11[m127 + b127*16 + a4*28*16] = data_11_array[a4][b127][m127];
        end
    endgenerate
    generate 
        localparam integer b128 = 16;
        for (m128 = 0; m128 < 16; m128 = m128 + 1) 
        begin: inbit128
            assign data_11[m128 + b128*16 + a4*28*16] = data_11_array[a4][b128][m128];
        end
    endgenerate
    generate 
        localparam integer b129 = 17;
        for (m129 = 0; m129 < 16; m129 = m129 + 1) 
        begin: inbit129
            assign data_11[m129 + b129*16 + a4*28*16] = data_11_array[a4][b129][m129];
        end
    endgenerate
    generate 
        localparam integer b130 = 18;
        for (m130 = 0; m130 < 16; m130 = m130 + 1) 
        begin: inbit130
            assign data_11[m130 + b130*16 + a4*28*16] = data_11_array[a4][b130][m130];
        end
    endgenerate
    generate 
        localparam integer b131 = 19;
        for (m131 = 0; m131 < 16; m131 = m131 + 1) 
        begin: inbit131
            assign data_11[m131 + b131*16 + a4*28*16] = data_11_array[a4][b131][m131];
        end
    endgenerate
    generate 
        localparam integer b132 = 20;
        for (m132 = 0; m132 < 16; m132 = m132 + 1) 
        begin: inbit132
            assign data_11[m132 + b132*16 + a4*28*16] = data_11_array[a4][b132][m132];
        end
    endgenerate
    generate 
        localparam integer b133 = 21;
        for (m133 = 0; m133 < 16; m133 = m133 + 1) 
        begin: inbit133
            assign data_11[m133 + b133*16 + a4*28*16] = data_11_array[a4][b133][m133];
        end
    endgenerate
    generate 
        localparam integer b134 = 22;
        for (m134 = 0; m134 < 16; m134 = m134 + 1) 
        begin: inbit134
            assign data_11[m134 + b134*16 + a4*28*16] = data_11_array[a4][b134][m134];
        end
    endgenerate
    generate 
        localparam integer b135 = 23;
        for (m135 = 0; m135 < 16; m135 = m135 + 1) 
        begin: inbit135
            assign data_11[m135 + b135*16 + a4*28*16] = data_11_array[a4][b135][m135];
        end
    endgenerate
    generate 
        localparam integer b136 = 24;
        for (m136 = 0; m136 < 16; m136 = m136 + 1) 
        begin: inbit136
            assign data_11[m136 + b136*16 + a4*28*16] = data_11_array[a4][b136][m136];
        end
    endgenerate
    generate 
        localparam integer b137 = 25;
        for (m137 = 0; m137 < 16; m137 = m137 + 1) 
        begin: inbit137
            assign data_11[m137 + b137*16 + a4*28*16] = data_11_array[a4][b137][m137];
        end
    endgenerate
    generate 
        localparam integer b138 = 26;
        for (m138 = 0; m138 < 16; m138 = m138 + 1) 
        begin: inbit138
            assign data_11[m138 + b138*16 + a4*28*16] = data_11_array[a4][b138][m138];
        end
    endgenerate
    generate 
        localparam integer b139 = 27;
        for (m139 = 0; m139 < 16; m139 = m139 + 1) 
        begin: inbit139
            assign data_11[m139 + b139*16 + a4*28*16] = data_11_array[a4][b139][m139];
        end
    endgenerate
    localparam integer a5 = 5;
    generate 
        localparam integer b140 = 0;
        for (m140 = 0; m140 < 16; m140 = m140 + 1) 
        begin: inbit140
            assign data_11[m140 + b140*16 + a5*28*16] = data_11_array[a5][b140][m140];
        end
    endgenerate
    generate 
        localparam integer b141 = 1;
        for (m141 = 0; m141 < 16; m141 = m141 + 1) 
        begin: inbit141
            assign data_11[m141 + b141*16 + a5*28*16] = data_11_array[a5][b141][m141];
        end
    endgenerate
    generate 
        localparam integer b142 = 2;
        for (m142 = 0; m142 < 16; m142 = m142 + 1) 
        begin: inbit142
            assign data_11[m142 + b142*16 + a5*28*16] = data_11_array[a5][b142][m142];
        end
    endgenerate
    generate 
        localparam integer b143 = 3;
        for (m143 = 0; m143 < 16; m143 = m143 + 1) 
        begin: inbit143
            assign data_11[m143 + b143*16 + a5*28*16] = data_11_array[a5][b143][m143];
        end
    endgenerate
    generate 
        localparam integer b144 = 4;
        for (m144 = 0; m144 < 16; m144 = m144 + 1) 
        begin: inbit144
            assign data_11[m144 + b144*16 + a5*28*16] = data_11_array[a5][b144][m144];
        end
    endgenerate
    generate 
        localparam integer b145 = 5;
        for (m145 = 0; m145 < 16; m145 = m145 + 1) 
        begin: inbit145
            assign data_11[m145 + b145*16 + a5*28*16] = data_11_array[a5][b145][m145];
        end
    endgenerate
    generate 
        localparam integer b146 = 6;
        for (m146 = 0; m146 < 16; m146 = m146 + 1) 
        begin: inbit146
            assign data_11[m146 + b146*16 + a5*28*16] = data_11_array[a5][b146][m146];
        end
    endgenerate
    generate 
        localparam integer b147 = 7;
        for (m147 = 0; m147 < 16; m147 = m147 + 1) 
        begin: inbit147
            assign data_11[m147 + b147*16 + a5*28*16] = data_11_array[a5][b147][m147];
        end
    endgenerate
    generate 
        localparam integer b148 = 8;
        for (m148 = 0; m148 < 16; m148 = m148 + 1) 
        begin: inbit148
            assign data_11[m148 + b148*16 + a5*28*16] = data_11_array[a5][b148][m148];
        end
    endgenerate
    generate 
        localparam integer b149 = 9;
        for (m149 = 0; m149 < 16; m149 = m149 + 1) 
        begin: inbit149
            assign data_11[m149 + b149*16 + a5*28*16] = data_11_array[a5][b149][m149];
        end
    endgenerate
    generate 
        localparam integer b150 = 10;
        for (m150 = 0; m150 < 16; m150 = m150 + 1) 
        begin: inbit150
            assign data_11[m150 + b150*16 + a5*28*16] = data_11_array[a5][b150][m150];
        end
    endgenerate
    generate 
        localparam integer b151 = 11;
        for (m151 = 0; m151 < 16; m151 = m151 + 1) 
        begin: inbit151
            assign data_11[m151 + b151*16 + a5*28*16] = data_11_array[a5][b151][m151];
        end
    endgenerate
    generate 
        localparam integer b152 = 12;
        for (m152 = 0; m152 < 16; m152 = m152 + 1) 
        begin: inbit152
            assign data_11[m152 + b152*16 + a5*28*16] = data_11_array[a5][b152][m152];
        end
    endgenerate
    generate 
        localparam integer b153 = 13;
        for (m153 = 0; m153 < 16; m153 = m153 + 1) 
        begin: inbit153
            assign data_11[m153 + b153*16 + a5*28*16] = data_11_array[a5][b153][m153];
        end
    endgenerate
    generate 
        localparam integer b154 = 14;
        for (m154 = 0; m154 < 16; m154 = m154 + 1) 
        begin: inbit154
            assign data_11[m154 + b154*16 + a5*28*16] = data_11_array[a5][b154][m154];
        end
    endgenerate
    generate 
        localparam integer b155 = 15;
        for (m155 = 0; m155 < 16; m155 = m155 + 1) 
        begin: inbit155
            assign data_11[m155 + b155*16 + a5*28*16] = data_11_array[a5][b155][m155];
        end
    endgenerate
    generate 
        localparam integer b156 = 16;
        for (m156 = 0; m156 < 16; m156 = m156 + 1) 
        begin: inbit156
            assign data_11[m156 + b156*16 + a5*28*16] = data_11_array[a5][b156][m156];
        end
    endgenerate
    generate 
        localparam integer b157 = 17;
        for (m157 = 0; m157 < 16; m157 = m157 + 1) 
        begin: inbit157
            assign data_11[m157 + b157*16 + a5*28*16] = data_11_array[a5][b157][m157];
        end
    endgenerate
    generate 
        localparam integer b158 = 18;
        for (m158 = 0; m158 < 16; m158 = m158 + 1) 
        begin: inbit158
            assign data_11[m158 + b158*16 + a5*28*16] = data_11_array[a5][b158][m158];
        end
    endgenerate
    generate 
        localparam integer b159 = 19;
        for (m159 = 0; m159 < 16; m159 = m159 + 1) 
        begin: inbit159
            assign data_11[m159 + b159*16 + a5*28*16] = data_11_array[a5][b159][m159];
        end
    endgenerate
    generate 
        localparam integer b160 = 20;
        for (m160 = 0; m160 < 16; m160 = m160 + 1) 
        begin: inbit160
            assign data_11[m160 + b160*16 + a5*28*16] = data_11_array[a5][b160][m160];
        end
    endgenerate
    generate 
        localparam integer b161 = 21;
        for (m161 = 0; m161 < 16; m161 = m161 + 1) 
        begin: inbit161
            assign data_11[m161 + b161*16 + a5*28*16] = data_11_array[a5][b161][m161];
        end
    endgenerate
    generate 
        localparam integer b162 = 22;
        for (m162 = 0; m162 < 16; m162 = m162 + 1) 
        begin: inbit162
            assign data_11[m162 + b162*16 + a5*28*16] = data_11_array[a5][b162][m162];
        end
    endgenerate
    generate 
        localparam integer b163 = 23;
        for (m163 = 0; m163 < 16; m163 = m163 + 1) 
        begin: inbit163
            assign data_11[m163 + b163*16 + a5*28*16] = data_11_array[a5][b163][m163];
        end
    endgenerate
    generate 
        localparam integer b164 = 24;
        for (m164 = 0; m164 < 16; m164 = m164 + 1) 
        begin: inbit164
            assign data_11[m164 + b164*16 + a5*28*16] = data_11_array[a5][b164][m164];
        end
    endgenerate
    generate 
        localparam integer b165 = 25;
        for (m165 = 0; m165 < 16; m165 = m165 + 1) 
        begin: inbit165
            assign data_11[m165 + b165*16 + a5*28*16] = data_11_array[a5][b165][m165];
        end
    endgenerate
    generate 
        localparam integer b166 = 26;
        for (m166 = 0; m166 < 16; m166 = m166 + 1) 
        begin: inbit166
            assign data_11[m166 + b166*16 + a5*28*16] = data_11_array[a5][b166][m166];
        end
    endgenerate
    generate 
        localparam integer b167 = 27;
        for (m167 = 0; m167 < 16; m167 = m167 + 1) 
        begin: inbit167
            assign data_11[m167 + b167*16 + a5*28*16] = data_11_array[a5][b167][m167];
        end
    endgenerate
    localparam integer a6 = 6;
    generate 
        localparam integer b168 = 0;
        for (m168 = 0; m168 < 16; m168 = m168 + 1) 
        begin: inbit168
            assign data_11[m168 + b168*16 + a6*28*16] = data_11_array[a6][b168][m168];
        end
    endgenerate
    generate 
        localparam integer b169 = 1;
        for (m169 = 0; m169 < 16; m169 = m169 + 1) 
        begin: inbit169
            assign data_11[m169 + b169*16 + a6*28*16] = data_11_array[a6][b169][m169];
        end
    endgenerate
    generate 
        localparam integer b170 = 2;
        for (m170 = 0; m170 < 16; m170 = m170 + 1) 
        begin: inbit170
            assign data_11[m170 + b170*16 + a6*28*16] = data_11_array[a6][b170][m170];
        end
    endgenerate
    generate 
        localparam integer b171 = 3;
        for (m171 = 0; m171 < 16; m171 = m171 + 1) 
        begin: inbit171
            assign data_11[m171 + b171*16 + a6*28*16] = data_11_array[a6][b171][m171];
        end
    endgenerate
    generate 
        localparam integer b172 = 4;
        for (m172 = 0; m172 < 16; m172 = m172 + 1) 
        begin: inbit172
            assign data_11[m172 + b172*16 + a6*28*16] = data_11_array[a6][b172][m172];
        end
    endgenerate
    generate 
        localparam integer b173 = 5;
        for (m173 = 0; m173 < 16; m173 = m173 + 1) 
        begin: inbit173
            assign data_11[m173 + b173*16 + a6*28*16] = data_11_array[a6][b173][m173];
        end
    endgenerate
    generate 
        localparam integer b174 = 6;
        for (m174 = 0; m174 < 16; m174 = m174 + 1) 
        begin: inbit174
            assign data_11[m174 + b174*16 + a6*28*16] = data_11_array[a6][b174][m174];
        end
    endgenerate
    generate 
        localparam integer b175 = 7;
        for (m175 = 0; m175 < 16; m175 = m175 + 1) 
        begin: inbit175
            assign data_11[m175 + b175*16 + a6*28*16] = data_11_array[a6][b175][m175];
        end
    endgenerate
    generate 
        localparam integer b176 = 8;
        for (m176 = 0; m176 < 16; m176 = m176 + 1) 
        begin: inbit176
            assign data_11[m176 + b176*16 + a6*28*16] = data_11_array[a6][b176][m176];
        end
    endgenerate
    generate 
        localparam integer b177 = 9;
        for (m177 = 0; m177 < 16; m177 = m177 + 1) 
        begin: inbit177
            assign data_11[m177 + b177*16 + a6*28*16] = data_11_array[a6][b177][m177];
        end
    endgenerate
    generate 
        localparam integer b178 = 10;
        for (m178 = 0; m178 < 16; m178 = m178 + 1) 
        begin: inbit178
            assign data_11[m178 + b178*16 + a6*28*16] = data_11_array[a6][b178][m178];
        end
    endgenerate
    generate 
        localparam integer b179 = 11;
        for (m179 = 0; m179 < 16; m179 = m179 + 1) 
        begin: inbit179
            assign data_11[m179 + b179*16 + a6*28*16] = data_11_array[a6][b179][m179];
        end
    endgenerate
    generate 
        localparam integer b180 = 12;
        for (m180 = 0; m180 < 16; m180 = m180 + 1) 
        begin: inbit180
            assign data_11[m180 + b180*16 + a6*28*16] = data_11_array[a6][b180][m180];
        end
    endgenerate
    generate 
        localparam integer b181 = 13;
        for (m181 = 0; m181 < 16; m181 = m181 + 1) 
        begin: inbit181
            assign data_11[m181 + b181*16 + a6*28*16] = data_11_array[a6][b181][m181];
        end
    endgenerate
    generate 
        localparam integer b182 = 14;
        for (m182 = 0; m182 < 16; m182 = m182 + 1) 
        begin: inbit182
            assign data_11[m182 + b182*16 + a6*28*16] = data_11_array[a6][b182][m182];
        end
    endgenerate
    generate 
        localparam integer b183 = 15;
        for (m183 = 0; m183 < 16; m183 = m183 + 1) 
        begin: inbit183
            assign data_11[m183 + b183*16 + a6*28*16] = data_11_array[a6][b183][m183];
        end
    endgenerate
    generate 
        localparam integer b184 = 16;
        for (m184 = 0; m184 < 16; m184 = m184 + 1) 
        begin: inbit184
            assign data_11[m184 + b184*16 + a6*28*16] = data_11_array[a6][b184][m184];
        end
    endgenerate
    generate 
        localparam integer b185 = 17;
        for (m185 = 0; m185 < 16; m185 = m185 + 1) 
        begin: inbit185
            assign data_11[m185 + b185*16 + a6*28*16] = data_11_array[a6][b185][m185];
        end
    endgenerate
    generate 
        localparam integer b186 = 18;
        for (m186 = 0; m186 < 16; m186 = m186 + 1) 
        begin: inbit186
            assign data_11[m186 + b186*16 + a6*28*16] = data_11_array[a6][b186][m186];
        end
    endgenerate
    generate 
        localparam integer b187 = 19;
        for (m187 = 0; m187 < 16; m187 = m187 + 1) 
        begin: inbit187
            assign data_11[m187 + b187*16 + a6*28*16] = data_11_array[a6][b187][m187];
        end
    endgenerate
    generate 
        localparam integer b188 = 20;
        for (m188 = 0; m188 < 16; m188 = m188 + 1) 
        begin: inbit188
            assign data_11[m188 + b188*16 + a6*28*16] = data_11_array[a6][b188][m188];
        end
    endgenerate
    generate 
        localparam integer b189 = 21;
        for (m189 = 0; m189 < 16; m189 = m189 + 1) 
        begin: inbit189
            assign data_11[m189 + b189*16 + a6*28*16] = data_11_array[a6][b189][m189];
        end
    endgenerate
    generate 
        localparam integer b190 = 22;
        for (m190 = 0; m190 < 16; m190 = m190 + 1) 
        begin: inbit190
            assign data_11[m190 + b190*16 + a6*28*16] = data_11_array[a6][b190][m190];
        end
    endgenerate
    generate 
        localparam integer b191 = 23;
        for (m191 = 0; m191 < 16; m191 = m191 + 1) 
        begin: inbit191
            assign data_11[m191 + b191*16 + a6*28*16] = data_11_array[a6][b191][m191];
        end
    endgenerate
    generate 
        localparam integer b192 = 24;
        for (m192 = 0; m192 < 16; m192 = m192 + 1) 
        begin: inbit192
            assign data_11[m192 + b192*16 + a6*28*16] = data_11_array[a6][b192][m192];
        end
    endgenerate
    generate 
        localparam integer b193 = 25;
        for (m193 = 0; m193 < 16; m193 = m193 + 1) 
        begin: inbit193
            assign data_11[m193 + b193*16 + a6*28*16] = data_11_array[a6][b193][m193];
        end
    endgenerate
    generate 
        localparam integer b194 = 26;
        for (m194 = 0; m194 < 16; m194 = m194 + 1) 
        begin: inbit194
            assign data_11[m194 + b194*16 + a6*28*16] = data_11_array[a6][b194][m194];
        end
    endgenerate
    generate 
        localparam integer b195 = 27;
        for (m195 = 0; m195 < 16; m195 = m195 + 1) 
        begin: inbit195
            assign data_11[m195 + b195*16 + a6*28*16] = data_11_array[a6][b195][m195];
        end
    endgenerate
    localparam integer a7 = 7;
    generate 
        localparam integer b196 = 0;
        for (m196 = 0; m196 < 16; m196 = m196 + 1) 
        begin: inbit196
            assign data_11[m196 + b196*16 + a7*28*16] = data_11_array[a7][b196][m196];
        end
    endgenerate
    generate 
        localparam integer b197 = 1;
        for (m197 = 0; m197 < 16; m197 = m197 + 1) 
        begin: inbit197
            assign data_11[m197 + b197*16 + a7*28*16] = data_11_array[a7][b197][m197];
        end
    endgenerate
    generate 
        localparam integer b198 = 2;
        for (m198 = 0; m198 < 16; m198 = m198 + 1) 
        begin: inbit198
            assign data_11[m198 + b198*16 + a7*28*16] = data_11_array[a7][b198][m198];
        end
    endgenerate
    generate 
        localparam integer b199 = 3;
        for (m199 = 0; m199 < 16; m199 = m199 + 1) 
        begin: inbit199
            assign data_11[m199 + b199*16 + a7*28*16] = data_11_array[a7][b199][m199];
        end
    endgenerate
    generate 
        localparam integer b200 = 4;
        for (m200 = 0; m200 < 16; m200 = m200 + 1) 
        begin: inbit200
            assign data_11[m200 + b200*16 + a7*28*16] = data_11_array[a7][b200][m200];
        end
    endgenerate
    generate 
        localparam integer b201 = 5;
        for (m201 = 0; m201 < 16; m201 = m201 + 1) 
        begin: inbit201
            assign data_11[m201 + b201*16 + a7*28*16] = data_11_array[a7][b201][m201];
        end
    endgenerate
    generate 
        localparam integer b202 = 6;
        for (m202 = 0; m202 < 16; m202 = m202 + 1) 
        begin: inbit202
            assign data_11[m202 + b202*16 + a7*28*16] = data_11_array[a7][b202][m202];
        end
    endgenerate
    generate 
        localparam integer b203 = 7;
        for (m203 = 0; m203 < 16; m203 = m203 + 1) 
        begin: inbit203
            assign data_11[m203 + b203*16 + a7*28*16] = data_11_array[a7][b203][m203];
        end
    endgenerate
    generate 
        localparam integer b204 = 8;
        for (m204 = 0; m204 < 16; m204 = m204 + 1) 
        begin: inbit204
            assign data_11[m204 + b204*16 + a7*28*16] = data_11_array[a7][b204][m204];
        end
    endgenerate
    generate 
        localparam integer b205 = 9;
        for (m205 = 0; m205 < 16; m205 = m205 + 1) 
        begin: inbit205
            assign data_11[m205 + b205*16 + a7*28*16] = data_11_array[a7][b205][m205];
        end
    endgenerate
    generate 
        localparam integer b206 = 10;
        for (m206 = 0; m206 < 16; m206 = m206 + 1) 
        begin: inbit206
            assign data_11[m206 + b206*16 + a7*28*16] = data_11_array[a7][b206][m206];
        end
    endgenerate
    generate 
        localparam integer b207 = 11;
        for (m207 = 0; m207 < 16; m207 = m207 + 1) 
        begin: inbit207
            assign data_11[m207 + b207*16 + a7*28*16] = data_11_array[a7][b207][m207];
        end
    endgenerate
    generate 
        localparam integer b208 = 12;
        for (m208 = 0; m208 < 16; m208 = m208 + 1) 
        begin: inbit208
            assign data_11[m208 + b208*16 + a7*28*16] = data_11_array[a7][b208][m208];
        end
    endgenerate
    generate 
        localparam integer b209 = 13;
        for (m209 = 0; m209 < 16; m209 = m209 + 1) 
        begin: inbit209
            assign data_11[m209 + b209*16 + a7*28*16] = data_11_array[a7][b209][m209];
        end
    endgenerate
    generate 
        localparam integer b210 = 14;
        for (m210 = 0; m210 < 16; m210 = m210 + 1) 
        begin: inbit210
            assign data_11[m210 + b210*16 + a7*28*16] = data_11_array[a7][b210][m210];
        end
    endgenerate
    generate 
        localparam integer b211 = 15;
        for (m211 = 0; m211 < 16; m211 = m211 + 1) 
        begin: inbit211
            assign data_11[m211 + b211*16 + a7*28*16] = data_11_array[a7][b211][m211];
        end
    endgenerate
    generate 
        localparam integer b212 = 16;
        for (m212 = 0; m212 < 16; m212 = m212 + 1) 
        begin: inbit212
            assign data_11[m212 + b212*16 + a7*28*16] = data_11_array[a7][b212][m212];
        end
    endgenerate
    generate 
        localparam integer b213 = 17;
        for (m213 = 0; m213 < 16; m213 = m213 + 1) 
        begin: inbit213
            assign data_11[m213 + b213*16 + a7*28*16] = data_11_array[a7][b213][m213];
        end
    endgenerate
    generate 
        localparam integer b214 = 18;
        for (m214 = 0; m214 < 16; m214 = m214 + 1) 
        begin: inbit214
            assign data_11[m214 + b214*16 + a7*28*16] = data_11_array[a7][b214][m214];
        end
    endgenerate
    generate 
        localparam integer b215 = 19;
        for (m215 = 0; m215 < 16; m215 = m215 + 1) 
        begin: inbit215
            assign data_11[m215 + b215*16 + a7*28*16] = data_11_array[a7][b215][m215];
        end
    endgenerate
    generate 
        localparam integer b216 = 20;
        for (m216 = 0; m216 < 16; m216 = m216 + 1) 
        begin: inbit216
            assign data_11[m216 + b216*16 + a7*28*16] = data_11_array[a7][b216][m216];
        end
    endgenerate
    generate 
        localparam integer b217 = 21;
        for (m217 = 0; m217 < 16; m217 = m217 + 1) 
        begin: inbit217
            assign data_11[m217 + b217*16 + a7*28*16] = data_11_array[a7][b217][m217];
        end
    endgenerate
    generate 
        localparam integer b218 = 22;
        for (m218 = 0; m218 < 16; m218 = m218 + 1) 
        begin: inbit218
            assign data_11[m218 + b218*16 + a7*28*16] = data_11_array[a7][b218][m218];
        end
    endgenerate
    generate 
        localparam integer b219 = 23;
        for (m219 = 0; m219 < 16; m219 = m219 + 1) 
        begin: inbit219
            assign data_11[m219 + b219*16 + a7*28*16] = data_11_array[a7][b219][m219];
        end
    endgenerate
    generate 
        localparam integer b220 = 24;
        for (m220 = 0; m220 < 16; m220 = m220 + 1) 
        begin: inbit220
            assign data_11[m220 + b220*16 + a7*28*16] = data_11_array[a7][b220][m220];
        end
    endgenerate
    generate 
        localparam integer b221 = 25;
        for (m221 = 0; m221 < 16; m221 = m221 + 1) 
        begin: inbit221
            assign data_11[m221 + b221*16 + a7*28*16] = data_11_array[a7][b221][m221];
        end
    endgenerate
    generate 
        localparam integer b222 = 26;
        for (m222 = 0; m222 < 16; m222 = m222 + 1) 
        begin: inbit222
            assign data_11[m222 + b222*16 + a7*28*16] = data_11_array[a7][b222][m222];
        end
    endgenerate
    generate 
        localparam integer b223 = 27;
        for (m223 = 0; m223 < 16; m223 = m223 + 1) 
        begin: inbit223
            assign data_11[m223 + b223*16 + a7*28*16] = data_11_array[a7][b223][m223];
        end
    endgenerate
    localparam integer a8 = 8;
    generate 
        localparam integer b224 = 0;
        for (m224 = 0; m224 < 16; m224 = m224 + 1) 
        begin: inbit224
            assign data_11[m224 + b224*16 + a8*28*16] = data_11_array[a8][b224][m224];
        end
    endgenerate
    generate 
        localparam integer b225 = 1;
        for (m225 = 0; m225 < 16; m225 = m225 + 1) 
        begin: inbit225
            assign data_11[m225 + b225*16 + a8*28*16] = data_11_array[a8][b225][m225];
        end
    endgenerate
    generate 
        localparam integer b226 = 2;
        for (m226 = 0; m226 < 16; m226 = m226 + 1) 
        begin: inbit226
            assign data_11[m226 + b226*16 + a8*28*16] = data_11_array[a8][b226][m226];
        end
    endgenerate
    generate 
        localparam integer b227 = 3;
        for (m227 = 0; m227 < 16; m227 = m227 + 1) 
        begin: inbit227
            assign data_11[m227 + b227*16 + a8*28*16] = data_11_array[a8][b227][m227];
        end
    endgenerate
    generate 
        localparam integer b228 = 4;
        for (m228 = 0; m228 < 16; m228 = m228 + 1) 
        begin: inbit228
            assign data_11[m228 + b228*16 + a8*28*16] = data_11_array[a8][b228][m228];
        end
    endgenerate
    generate 
        localparam integer b229 = 5;
        for (m229 = 0; m229 < 16; m229 = m229 + 1) 
        begin: inbit229
            assign data_11[m229 + b229*16 + a8*28*16] = data_11_array[a8][b229][m229];
        end
    endgenerate
    generate 
        localparam integer b230 = 6;
        for (m230 = 0; m230 < 16; m230 = m230 + 1) 
        begin: inbit230
            assign data_11[m230 + b230*16 + a8*28*16] = data_11_array[a8][b230][m230];
        end
    endgenerate
    generate 
        localparam integer b231 = 7;
        for (m231 = 0; m231 < 16; m231 = m231 + 1) 
        begin: inbit231
            assign data_11[m231 + b231*16 + a8*28*16] = data_11_array[a8][b231][m231];
        end
    endgenerate
    generate 
        localparam integer b232 = 8;
        for (m232 = 0; m232 < 16; m232 = m232 + 1) 
        begin: inbit232
            assign data_11[m232 + b232*16 + a8*28*16] = data_11_array[a8][b232][m232];
        end
    endgenerate
    generate 
        localparam integer b233 = 9;
        for (m233 = 0; m233 < 16; m233 = m233 + 1) 
        begin: inbit233
            assign data_11[m233 + b233*16 + a8*28*16] = data_11_array[a8][b233][m233];
        end
    endgenerate
    generate 
        localparam integer b234 = 10;
        for (m234 = 0; m234 < 16; m234 = m234 + 1) 
        begin: inbit234
            assign data_11[m234 + b234*16 + a8*28*16] = data_11_array[a8][b234][m234];
        end
    endgenerate
    generate 
        localparam integer b235 = 11;
        for (m235 = 0; m235 < 16; m235 = m235 + 1) 
        begin: inbit235
            assign data_11[m235 + b235*16 + a8*28*16] = data_11_array[a8][b235][m235];
        end
    endgenerate
    generate 
        localparam integer b236 = 12;
        for (m236 = 0; m236 < 16; m236 = m236 + 1) 
        begin: inbit236
            assign data_11[m236 + b236*16 + a8*28*16] = data_11_array[a8][b236][m236];
        end
    endgenerate
    generate 
        localparam integer b237 = 13;
        for (m237 = 0; m237 < 16; m237 = m237 + 1) 
        begin: inbit237
            assign data_11[m237 + b237*16 + a8*28*16] = data_11_array[a8][b237][m237];
        end
    endgenerate
    generate 
        localparam integer b238 = 14;
        for (m238 = 0; m238 < 16; m238 = m238 + 1) 
        begin: inbit238
            assign data_11[m238 + b238*16 + a8*28*16] = data_11_array[a8][b238][m238];
        end
    endgenerate
    generate 
        localparam integer b239 = 15;
        for (m239 = 0; m239 < 16; m239 = m239 + 1) 
        begin: inbit239
            assign data_11[m239 + b239*16 + a8*28*16] = data_11_array[a8][b239][m239];
        end
    endgenerate
    generate 
        localparam integer b240 = 16;
        for (m240 = 0; m240 < 16; m240 = m240 + 1) 
        begin: inbit240
            assign data_11[m240 + b240*16 + a8*28*16] = data_11_array[a8][b240][m240];
        end
    endgenerate
    generate 
        localparam integer b241 = 17;
        for (m241 = 0; m241 < 16; m241 = m241 + 1) 
        begin: inbit241
            assign data_11[m241 + b241*16 + a8*28*16] = data_11_array[a8][b241][m241];
        end
    endgenerate
    generate 
        localparam integer b242 = 18;
        for (m242 = 0; m242 < 16; m242 = m242 + 1) 
        begin: inbit242
            assign data_11[m242 + b242*16 + a8*28*16] = data_11_array[a8][b242][m242];
        end
    endgenerate
    generate 
        localparam integer b243 = 19;
        for (m243 = 0; m243 < 16; m243 = m243 + 1) 
        begin: inbit243
            assign data_11[m243 + b243*16 + a8*28*16] = data_11_array[a8][b243][m243];
        end
    endgenerate
    generate 
        localparam integer b244 = 20;
        for (m244 = 0; m244 < 16; m244 = m244 + 1) 
        begin: inbit244
            assign data_11[m244 + b244*16 + a8*28*16] = data_11_array[a8][b244][m244];
        end
    endgenerate
    generate 
        localparam integer b245 = 21;
        for (m245 = 0; m245 < 16; m245 = m245 + 1) 
        begin: inbit245
            assign data_11[m245 + b245*16 + a8*28*16] = data_11_array[a8][b245][m245];
        end
    endgenerate
    generate 
        localparam integer b246 = 22;
        for (m246 = 0; m246 < 16; m246 = m246 + 1) 
        begin: inbit246
            assign data_11[m246 + b246*16 + a8*28*16] = data_11_array[a8][b246][m246];
        end
    endgenerate
    generate 
        localparam integer b247 = 23;
        for (m247 = 0; m247 < 16; m247 = m247 + 1) 
        begin: inbit247
            assign data_11[m247 + b247*16 + a8*28*16] = data_11_array[a8][b247][m247];
        end
    endgenerate
    generate 
        localparam integer b248 = 24;
        for (m248 = 0; m248 < 16; m248 = m248 + 1) 
        begin: inbit248
            assign data_11[m248 + b248*16 + a8*28*16] = data_11_array[a8][b248][m248];
        end
    endgenerate
    generate 
        localparam integer b249 = 25;
        for (m249 = 0; m249 < 16; m249 = m249 + 1) 
        begin: inbit249
            assign data_11[m249 + b249*16 + a8*28*16] = data_11_array[a8][b249][m249];
        end
    endgenerate
    generate 
        localparam integer b250 = 26;
        for (m250 = 0; m250 < 16; m250 = m250 + 1) 
        begin: inbit250
            assign data_11[m250 + b250*16 + a8*28*16] = data_11_array[a8][b250][m250];
        end
    endgenerate
    generate 
        localparam integer b251 = 27;
        for (m251 = 0; m251 < 16; m251 = m251 + 1) 
        begin: inbit251
            assign data_11[m251 + b251*16 + a8*28*16] = data_11_array[a8][b251][m251];
        end
    endgenerate
    localparam integer a9 = 9;
    generate 
        localparam integer b252 = 0;
        for (m252 = 0; m252 < 16; m252 = m252 + 1) 
        begin: inbit252
            assign data_11[m252 + b252*16 + a9*28*16] = data_11_array[a9][b252][m252];
        end
    endgenerate
    generate 
        localparam integer b253 = 1;
        for (m253 = 0; m253 < 16; m253 = m253 + 1) 
        begin: inbit253
            assign data_11[m253 + b253*16 + a9*28*16] = data_11_array[a9][b253][m253];
        end
    endgenerate
    generate 
        localparam integer b254 = 2;
        for (m254 = 0; m254 < 16; m254 = m254 + 1) 
        begin: inbit254
            assign data_11[m254 + b254*16 + a9*28*16] = data_11_array[a9][b254][m254];
        end
    endgenerate
    generate 
        localparam integer b255 = 3;
        for (m255 = 0; m255 < 16; m255 = m255 + 1) 
        begin: inbit255
            assign data_11[m255 + b255*16 + a9*28*16] = data_11_array[a9][b255][m255];
        end
    endgenerate
    generate 
        localparam integer b256 = 4;
        for (m256 = 0; m256 < 16; m256 = m256 + 1) 
        begin: inbit256
            assign data_11[m256 + b256*16 + a9*28*16] = data_11_array[a9][b256][m256];
        end
    endgenerate
    generate 
        localparam integer b257 = 5;
        for (m257 = 0; m257 < 16; m257 = m257 + 1) 
        begin: inbit257
            assign data_11[m257 + b257*16 + a9*28*16] = data_11_array[a9][b257][m257];
        end
    endgenerate
    generate 
        localparam integer b258 = 6;
        for (m258 = 0; m258 < 16; m258 = m258 + 1) 
        begin: inbit258
            assign data_11[m258 + b258*16 + a9*28*16] = data_11_array[a9][b258][m258];
        end
    endgenerate
    generate 
        localparam integer b259 = 7;
        for (m259 = 0; m259 < 16; m259 = m259 + 1) 
        begin: inbit259
            assign data_11[m259 + b259*16 + a9*28*16] = data_11_array[a9][b259][m259];
        end
    endgenerate
    generate 
        localparam integer b260 = 8;
        for (m260 = 0; m260 < 16; m260 = m260 + 1) 
        begin: inbit260
            assign data_11[m260 + b260*16 + a9*28*16] = data_11_array[a9][b260][m260];
        end
    endgenerate
    generate 
        localparam integer b261 = 9;
        for (m261 = 0; m261 < 16; m261 = m261 + 1) 
        begin: inbit261
            assign data_11[m261 + b261*16 + a9*28*16] = data_11_array[a9][b261][m261];
        end
    endgenerate
    generate 
        localparam integer b262 = 10;
        for (m262 = 0; m262 < 16; m262 = m262 + 1) 
        begin: inbit262
            assign data_11[m262 + b262*16 + a9*28*16] = data_11_array[a9][b262][m262];
        end
    endgenerate
    generate 
        localparam integer b263 = 11;
        for (m263 = 0; m263 < 16; m263 = m263 + 1) 
        begin: inbit263
            assign data_11[m263 + b263*16 + a9*28*16] = data_11_array[a9][b263][m263];
        end
    endgenerate
    generate 
        localparam integer b264 = 12;
        for (m264 = 0; m264 < 16; m264 = m264 + 1) 
        begin: inbit264
            assign data_11[m264 + b264*16 + a9*28*16] = data_11_array[a9][b264][m264];
        end
    endgenerate
    generate 
        localparam integer b265 = 13;
        for (m265 = 0; m265 < 16; m265 = m265 + 1) 
        begin: inbit265
            assign data_11[m265 + b265*16 + a9*28*16] = data_11_array[a9][b265][m265];
        end
    endgenerate
    generate 
        localparam integer b266 = 14;
        for (m266 = 0; m266 < 16; m266 = m266 + 1) 
        begin: inbit266
            assign data_11[m266 + b266*16 + a9*28*16] = data_11_array[a9][b266][m266];
        end
    endgenerate
    generate 
        localparam integer b267 = 15;
        for (m267 = 0; m267 < 16; m267 = m267 + 1) 
        begin: inbit267
            assign data_11[m267 + b267*16 + a9*28*16] = data_11_array[a9][b267][m267];
        end
    endgenerate
    generate 
        localparam integer b268 = 16;
        for (m268 = 0; m268 < 16; m268 = m268 + 1) 
        begin: inbit268
            assign data_11[m268 + b268*16 + a9*28*16] = data_11_array[a9][b268][m268];
        end
    endgenerate
    generate 
        localparam integer b269 = 17;
        for (m269 = 0; m269 < 16; m269 = m269 + 1) 
        begin: inbit269
            assign data_11[m269 + b269*16 + a9*28*16] = data_11_array[a9][b269][m269];
        end
    endgenerate
    generate 
        localparam integer b270 = 18;
        for (m270 = 0; m270 < 16; m270 = m270 + 1) 
        begin: inbit270
            assign data_11[m270 + b270*16 + a9*28*16] = data_11_array[a9][b270][m270];
        end
    endgenerate
    generate 
        localparam integer b271 = 19;
        for (m271 = 0; m271 < 16; m271 = m271 + 1) 
        begin: inbit271
            assign data_11[m271 + b271*16 + a9*28*16] = data_11_array[a9][b271][m271];
        end
    endgenerate
    generate 
        localparam integer b272 = 20;
        for (m272 = 0; m272 < 16; m272 = m272 + 1) 
        begin: inbit272
            assign data_11[m272 + b272*16 + a9*28*16] = data_11_array[a9][b272][m272];
        end
    endgenerate
    generate 
        localparam integer b273 = 21;
        for (m273 = 0; m273 < 16; m273 = m273 + 1) 
        begin: inbit273
            assign data_11[m273 + b273*16 + a9*28*16] = data_11_array[a9][b273][m273];
        end
    endgenerate
    generate 
        localparam integer b274 = 22;
        for (m274 = 0; m274 < 16; m274 = m274 + 1) 
        begin: inbit274
            assign data_11[m274 + b274*16 + a9*28*16] = data_11_array[a9][b274][m274];
        end
    endgenerate
    generate 
        localparam integer b275 = 23;
        for (m275 = 0; m275 < 16; m275 = m275 + 1) 
        begin: inbit275
            assign data_11[m275 + b275*16 + a9*28*16] = data_11_array[a9][b275][m275];
        end
    endgenerate
    generate 
        localparam integer b276 = 24;
        for (m276 = 0; m276 < 16; m276 = m276 + 1) 
        begin: inbit276
            assign data_11[m276 + b276*16 + a9*28*16] = data_11_array[a9][b276][m276];
        end
    endgenerate
    generate 
        localparam integer b277 = 25;
        for (m277 = 0; m277 < 16; m277 = m277 + 1) 
        begin: inbit277
            assign data_11[m277 + b277*16 + a9*28*16] = data_11_array[a9][b277][m277];
        end
    endgenerate
    generate 
        localparam integer b278 = 26;
        for (m278 = 0; m278 < 16; m278 = m278 + 1) 
        begin: inbit278
            assign data_11[m278 + b278*16 + a9*28*16] = data_11_array[a9][b278][m278];
        end
    endgenerate
    generate 
        localparam integer b279 = 27;
        for (m279 = 0; m279 < 16; m279 = m279 + 1) 
        begin: inbit279
            assign data_11[m279 + b279*16 + a9*28*16] = data_11_array[a9][b279][m279];
        end
    endgenerate
    localparam integer a10 = 10;
    generate 
        localparam integer b280 = 0;
        for (m280 = 0; m280 < 16; m280 = m280 + 1) 
        begin: inbit280
            assign data_11[m280 + b280*16 + a10*28*16] = data_11_array[a10][b280][m280];
        end
    endgenerate
    generate 
        localparam integer b281 = 1;
        for (m281 = 0; m281 < 16; m281 = m281 + 1) 
        begin: inbit281
            assign data_11[m281 + b281*16 + a10*28*16] = data_11_array[a10][b281][m281];
        end
    endgenerate
    generate 
        localparam integer b282 = 2;
        for (m282 = 0; m282 < 16; m282 = m282 + 1) 
        begin: inbit282
            assign data_11[m282 + b282*16 + a10*28*16] = data_11_array[a10][b282][m282];
        end
    endgenerate
    generate 
        localparam integer b283 = 3;
        for (m283 = 0; m283 < 16; m283 = m283 + 1) 
        begin: inbit283
            assign data_11[m283 + b283*16 + a10*28*16] = data_11_array[a10][b283][m283];
        end
    endgenerate
    generate 
        localparam integer b284 = 4;
        for (m284 = 0; m284 < 16; m284 = m284 + 1) 
        begin: inbit284
            assign data_11[m284 + b284*16 + a10*28*16] = data_11_array[a10][b284][m284];
        end
    endgenerate
    generate 
        localparam integer b285 = 5;
        for (m285 = 0; m285 < 16; m285 = m285 + 1) 
        begin: inbit285
            assign data_11[m285 + b285*16 + a10*28*16] = data_11_array[a10][b285][m285];
        end
    endgenerate
    generate 
        localparam integer b286 = 6;
        for (m286 = 0; m286 < 16; m286 = m286 + 1) 
        begin: inbit286
            assign data_11[m286 + b286*16 + a10*28*16] = data_11_array[a10][b286][m286];
        end
    endgenerate
    generate 
        localparam integer b287 = 7;
        for (m287 = 0; m287 < 16; m287 = m287 + 1) 
        begin: inbit287
            assign data_11[m287 + b287*16 + a10*28*16] = data_11_array[a10][b287][m287];
        end
    endgenerate
    generate 
        localparam integer b288 = 8;
        for (m288 = 0; m288 < 16; m288 = m288 + 1) 
        begin: inbit288
            assign data_11[m288 + b288*16 + a10*28*16] = data_11_array[a10][b288][m288];
        end
    endgenerate
    generate 
        localparam integer b289 = 9;
        for (m289 = 0; m289 < 16; m289 = m289 + 1) 
        begin: inbit289
            assign data_11[m289 + b289*16 + a10*28*16] = data_11_array[a10][b289][m289];
        end
    endgenerate
    generate 
        localparam integer b290 = 10;
        for (m290 = 0; m290 < 16; m290 = m290 + 1) 
        begin: inbit290
            assign data_11[m290 + b290*16 + a10*28*16] = data_11_array[a10][b290][m290];
        end
    endgenerate
    generate 
        localparam integer b291 = 11;
        for (m291 = 0; m291 < 16; m291 = m291 + 1) 
        begin: inbit291
            assign data_11[m291 + b291*16 + a10*28*16] = data_11_array[a10][b291][m291];
        end
    endgenerate
    generate 
        localparam integer b292 = 12;
        for (m292 = 0; m292 < 16; m292 = m292 + 1) 
        begin: inbit292
            assign data_11[m292 + b292*16 + a10*28*16] = data_11_array[a10][b292][m292];
        end
    endgenerate
    generate 
        localparam integer b293 = 13;
        for (m293 = 0; m293 < 16; m293 = m293 + 1) 
        begin: inbit293
            assign data_11[m293 + b293*16 + a10*28*16] = data_11_array[a10][b293][m293];
        end
    endgenerate
    generate 
        localparam integer b294 = 14;
        for (m294 = 0; m294 < 16; m294 = m294 + 1) 
        begin: inbit294
            assign data_11[m294 + b294*16 + a10*28*16] = data_11_array[a10][b294][m294];
        end
    endgenerate
    generate 
        localparam integer b295 = 15;
        for (m295 = 0; m295 < 16; m295 = m295 + 1) 
        begin: inbit295
            assign data_11[m295 + b295*16 + a10*28*16] = data_11_array[a10][b295][m295];
        end
    endgenerate
    generate 
        localparam integer b296 = 16;
        for (m296 = 0; m296 < 16; m296 = m296 + 1) 
        begin: inbit296
            assign data_11[m296 + b296*16 + a10*28*16] = data_11_array[a10][b296][m296];
        end
    endgenerate
    generate 
        localparam integer b297 = 17;
        for (m297 = 0; m297 < 16; m297 = m297 + 1) 
        begin: inbit297
            assign data_11[m297 + b297*16 + a10*28*16] = data_11_array[a10][b297][m297];
        end
    endgenerate
    generate 
        localparam integer b298 = 18;
        for (m298 = 0; m298 < 16; m298 = m298 + 1) 
        begin: inbit298
            assign data_11[m298 + b298*16 + a10*28*16] = data_11_array[a10][b298][m298];
        end
    endgenerate
    generate 
        localparam integer b299 = 19;
        for (m299 = 0; m299 < 16; m299 = m299 + 1) 
        begin: inbit299
            assign data_11[m299 + b299*16 + a10*28*16] = data_11_array[a10][b299][m299];
        end
    endgenerate
    generate 
        localparam integer b300 = 20;
        for (m300 = 0; m300 < 16; m300 = m300 + 1) 
        begin: inbit300
            assign data_11[m300 + b300*16 + a10*28*16] = data_11_array[a10][b300][m300];
        end
    endgenerate
    generate 
        localparam integer b301 = 21;
        for (m301 = 0; m301 < 16; m301 = m301 + 1) 
        begin: inbit301
            assign data_11[m301 + b301*16 + a10*28*16] = data_11_array[a10][b301][m301];
        end
    endgenerate
    generate 
        localparam integer b302 = 22;
        for (m302 = 0; m302 < 16; m302 = m302 + 1) 
        begin: inbit302
            assign data_11[m302 + b302*16 + a10*28*16] = data_11_array[a10][b302][m302];
        end
    endgenerate
    generate 
        localparam integer b303 = 23;
        for (m303 = 0; m303 < 16; m303 = m303 + 1) 
        begin: inbit303
            assign data_11[m303 + b303*16 + a10*28*16] = data_11_array[a10][b303][m303];
        end
    endgenerate
    generate 
        localparam integer b304 = 24;
        for (m304 = 0; m304 < 16; m304 = m304 + 1) 
        begin: inbit304
            assign data_11[m304 + b304*16 + a10*28*16] = data_11_array[a10][b304][m304];
        end
    endgenerate
    generate 
        localparam integer b305 = 25;
        for (m305 = 0; m305 < 16; m305 = m305 + 1) 
        begin: inbit305
            assign data_11[m305 + b305*16 + a10*28*16] = data_11_array[a10][b305][m305];
        end
    endgenerate
    generate 
        localparam integer b306 = 26;
        for (m306 = 0; m306 < 16; m306 = m306 + 1) 
        begin: inbit306
            assign data_11[m306 + b306*16 + a10*28*16] = data_11_array[a10][b306][m306];
        end
    endgenerate
    generate 
        localparam integer b307 = 27;
        for (m307 = 0; m307 < 16; m307 = m307 + 1) 
        begin: inbit307
            assign data_11[m307 + b307*16 + a10*28*16] = data_11_array[a10][b307][m307];
        end
    endgenerate
    localparam integer a11 = 11;
    generate 
        localparam integer b308 = 0;
        for (m308 = 0; m308 < 16; m308 = m308 + 1) 
        begin: inbit308
            assign data_11[m308 + b308*16 + a11*28*16] = data_11_array[a11][b308][m308];
        end
    endgenerate
    generate 
        localparam integer b309 = 1;
        for (m309 = 0; m309 < 16; m309 = m309 + 1) 
        begin: inbit309
            assign data_11[m309 + b309*16 + a11*28*16] = data_11_array[a11][b309][m309];
        end
    endgenerate
    generate 
        localparam integer b310 = 2;
        for (m310 = 0; m310 < 16; m310 = m310 + 1) 
        begin: inbit310
            assign data_11[m310 + b310*16 + a11*28*16] = data_11_array[a11][b310][m310];
        end
    endgenerate
    generate 
        localparam integer b311 = 3;
        for (m311 = 0; m311 < 16; m311 = m311 + 1) 
        begin: inbit311
            assign data_11[m311 + b311*16 + a11*28*16] = data_11_array[a11][b311][m311];
        end
    endgenerate
    generate 
        localparam integer b312 = 4;
        for (m312 = 0; m312 < 16; m312 = m312 + 1) 
        begin: inbit312
            assign data_11[m312 + b312*16 + a11*28*16] = data_11_array[a11][b312][m312];
        end
    endgenerate
    generate 
        localparam integer b313 = 5;
        for (m313 = 0; m313 < 16; m313 = m313 + 1) 
        begin: inbit313
            assign data_11[m313 + b313*16 + a11*28*16] = data_11_array[a11][b313][m313];
        end
    endgenerate
    generate 
        localparam integer b314 = 6;
        for (m314 = 0; m314 < 16; m314 = m314 + 1) 
        begin: inbit314
            assign data_11[m314 + b314*16 + a11*28*16] = data_11_array[a11][b314][m314];
        end
    endgenerate
    generate 
        localparam integer b315 = 7;
        for (m315 = 0; m315 < 16; m315 = m315 + 1) 
        begin: inbit315
            assign data_11[m315 + b315*16 + a11*28*16] = data_11_array[a11][b315][m315];
        end
    endgenerate
    generate 
        localparam integer b316 = 8;
        for (m316 = 0; m316 < 16; m316 = m316 + 1) 
        begin: inbit316
            assign data_11[m316 + b316*16 + a11*28*16] = data_11_array[a11][b316][m316];
        end
    endgenerate
    generate 
        localparam integer b317 = 9;
        for (m317 = 0; m317 < 16; m317 = m317 + 1) 
        begin: inbit317
            assign data_11[m317 + b317*16 + a11*28*16] = data_11_array[a11][b317][m317];
        end
    endgenerate
    generate 
        localparam integer b318 = 10;
        for (m318 = 0; m318 < 16; m318 = m318 + 1) 
        begin: inbit318
            assign data_11[m318 + b318*16 + a11*28*16] = data_11_array[a11][b318][m318];
        end
    endgenerate
    generate 
        localparam integer b319 = 11;
        for (m319 = 0; m319 < 16; m319 = m319 + 1) 
        begin: inbit319
            assign data_11[m319 + b319*16 + a11*28*16] = data_11_array[a11][b319][m319];
        end
    endgenerate
    generate 
        localparam integer b320 = 12;
        for (m320 = 0; m320 < 16; m320 = m320 + 1) 
        begin: inbit320
            assign data_11[m320 + b320*16 + a11*28*16] = data_11_array[a11][b320][m320];
        end
    endgenerate
    generate 
        localparam integer b321 = 13;
        for (m321 = 0; m321 < 16; m321 = m321 + 1) 
        begin: inbit321
            assign data_11[m321 + b321*16 + a11*28*16] = data_11_array[a11][b321][m321];
        end
    endgenerate
    generate 
        localparam integer b322 = 14;
        for (m322 = 0; m322 < 16; m322 = m322 + 1) 
        begin: inbit322
            assign data_11[m322 + b322*16 + a11*28*16] = data_11_array[a11][b322][m322];
        end
    endgenerate
    generate 
        localparam integer b323 = 15;
        for (m323 = 0; m323 < 16; m323 = m323 + 1) 
        begin: inbit323
            assign data_11[m323 + b323*16 + a11*28*16] = data_11_array[a11][b323][m323];
        end
    endgenerate
    generate 
        localparam integer b324 = 16;
        for (m324 = 0; m324 < 16; m324 = m324 + 1) 
        begin: inbit324
            assign data_11[m324 + b324*16 + a11*28*16] = data_11_array[a11][b324][m324];
        end
    endgenerate
    generate 
        localparam integer b325 = 17;
        for (m325 = 0; m325 < 16; m325 = m325 + 1) 
        begin: inbit325
            assign data_11[m325 + b325*16 + a11*28*16] = data_11_array[a11][b325][m325];
        end
    endgenerate
    generate 
        localparam integer b326 = 18;
        for (m326 = 0; m326 < 16; m326 = m326 + 1) 
        begin: inbit326
            assign data_11[m326 + b326*16 + a11*28*16] = data_11_array[a11][b326][m326];
        end
    endgenerate
    generate 
        localparam integer b327 = 19;
        for (m327 = 0; m327 < 16; m327 = m327 + 1) 
        begin: inbit327
            assign data_11[m327 + b327*16 + a11*28*16] = data_11_array[a11][b327][m327];
        end
    endgenerate
    generate 
        localparam integer b328 = 20;
        for (m328 = 0; m328 < 16; m328 = m328 + 1) 
        begin: inbit328
            assign data_11[m328 + b328*16 + a11*28*16] = data_11_array[a11][b328][m328];
        end
    endgenerate
    generate 
        localparam integer b329 = 21;
        for (m329 = 0; m329 < 16; m329 = m329 + 1) 
        begin: inbit329
            assign data_11[m329 + b329*16 + a11*28*16] = data_11_array[a11][b329][m329];
        end
    endgenerate
    generate 
        localparam integer b330 = 22;
        for (m330 = 0; m330 < 16; m330 = m330 + 1) 
        begin: inbit330
            assign data_11[m330 + b330*16 + a11*28*16] = data_11_array[a11][b330][m330];
        end
    endgenerate
    generate 
        localparam integer b331 = 23;
        for (m331 = 0; m331 < 16; m331 = m331 + 1) 
        begin: inbit331
            assign data_11[m331 + b331*16 + a11*28*16] = data_11_array[a11][b331][m331];
        end
    endgenerate
    generate 
        localparam integer b332 = 24;
        for (m332 = 0; m332 < 16; m332 = m332 + 1) 
        begin: inbit332
            assign data_11[m332 + b332*16 + a11*28*16] = data_11_array[a11][b332][m332];
        end
    endgenerate
    generate 
        localparam integer b333 = 25;
        for (m333 = 0; m333 < 16; m333 = m333 + 1) 
        begin: inbit333
            assign data_11[m333 + b333*16 + a11*28*16] = data_11_array[a11][b333][m333];
        end
    endgenerate
    generate 
        localparam integer b334 = 26;
        for (m334 = 0; m334 < 16; m334 = m334 + 1) 
        begin: inbit334
            assign data_11[m334 + b334*16 + a11*28*16] = data_11_array[a11][b334][m334];
        end
    endgenerate
    generate 
        localparam integer b335 = 27;
        for (m335 = 0; m335 < 16; m335 = m335 + 1) 
        begin: inbit335
            assign data_11[m335 + b335*16 + a11*28*16] = data_11_array[a11][b335][m335];
        end
    endgenerate
    localparam integer a12 = 12;
    generate 
        localparam integer b336 = 0;
        for (m336 = 0; m336 < 16; m336 = m336 + 1) 
        begin: inbit336
            assign data_11[m336 + b336*16 + a12*28*16] = data_11_array[a12][b336][m336];
        end
    endgenerate
    generate 
        localparam integer b337 = 1;
        for (m337 = 0; m337 < 16; m337 = m337 + 1) 
        begin: inbit337
            assign data_11[m337 + b337*16 + a12*28*16] = data_11_array[a12][b337][m337];
        end
    endgenerate
    generate 
        localparam integer b338 = 2;
        for (m338 = 0; m338 < 16; m338 = m338 + 1) 
        begin: inbit338
            assign data_11[m338 + b338*16 + a12*28*16] = data_11_array[a12][b338][m338];
        end
    endgenerate
    generate 
        localparam integer b339 = 3;
        for (m339 = 0; m339 < 16; m339 = m339 + 1) 
        begin: inbit339
            assign data_11[m339 + b339*16 + a12*28*16] = data_11_array[a12][b339][m339];
        end
    endgenerate
    generate 
        localparam integer b340 = 4;
        for (m340 = 0; m340 < 16; m340 = m340 + 1) 
        begin: inbit340
            assign data_11[m340 + b340*16 + a12*28*16] = data_11_array[a12][b340][m340];
        end
    endgenerate
    generate 
        localparam integer b341 = 5;
        for (m341 = 0; m341 < 16; m341 = m341 + 1) 
        begin: inbit341
            assign data_11[m341 + b341*16 + a12*28*16] = data_11_array[a12][b341][m341];
        end
    endgenerate
    generate 
        localparam integer b342 = 6;
        for (m342 = 0; m342 < 16; m342 = m342 + 1) 
        begin: inbit342
            assign data_11[m342 + b342*16 + a12*28*16] = data_11_array[a12][b342][m342];
        end
    endgenerate
    generate 
        localparam integer b343 = 7;
        for (m343 = 0; m343 < 16; m343 = m343 + 1) 
        begin: inbit343
            assign data_11[m343 + b343*16 + a12*28*16] = data_11_array[a12][b343][m343];
        end
    endgenerate
    generate 
        localparam integer b344 = 8;
        for (m344 = 0; m344 < 16; m344 = m344 + 1) 
        begin: inbit344
            assign data_11[m344 + b344*16 + a12*28*16] = data_11_array[a12][b344][m344];
        end
    endgenerate
    generate 
        localparam integer b345 = 9;
        for (m345 = 0; m345 < 16; m345 = m345 + 1) 
        begin: inbit345
            assign data_11[m345 + b345*16 + a12*28*16] = data_11_array[a12][b345][m345];
        end
    endgenerate
    generate 
        localparam integer b346 = 10;
        for (m346 = 0; m346 < 16; m346 = m346 + 1) 
        begin: inbit346
            assign data_11[m346 + b346*16 + a12*28*16] = data_11_array[a12][b346][m346];
        end
    endgenerate
    generate 
        localparam integer b347 = 11;
        for (m347 = 0; m347 < 16; m347 = m347 + 1) 
        begin: inbit347
            assign data_11[m347 + b347*16 + a12*28*16] = data_11_array[a12][b347][m347];
        end
    endgenerate
    generate 
        localparam integer b348 = 12;
        for (m348 = 0; m348 < 16; m348 = m348 + 1) 
        begin: inbit348
            assign data_11[m348 + b348*16 + a12*28*16] = data_11_array[a12][b348][m348];
        end
    endgenerate
    generate 
        localparam integer b349 = 13;
        for (m349 = 0; m349 < 16; m349 = m349 + 1) 
        begin: inbit349
            assign data_11[m349 + b349*16 + a12*28*16] = data_11_array[a12][b349][m349];
        end
    endgenerate
    generate 
        localparam integer b350 = 14;
        for (m350 = 0; m350 < 16; m350 = m350 + 1) 
        begin: inbit350
            assign data_11[m350 + b350*16 + a12*28*16] = data_11_array[a12][b350][m350];
        end
    endgenerate
    generate 
        localparam integer b351 = 15;
        for (m351 = 0; m351 < 16; m351 = m351 + 1) 
        begin: inbit351
            assign data_11[m351 + b351*16 + a12*28*16] = data_11_array[a12][b351][m351];
        end
    endgenerate
    generate 
        localparam integer b352 = 16;
        for (m352 = 0; m352 < 16; m352 = m352 + 1) 
        begin: inbit352
            assign data_11[m352 + b352*16 + a12*28*16] = data_11_array[a12][b352][m352];
        end
    endgenerate
    generate 
        localparam integer b353 = 17;
        for (m353 = 0; m353 < 16; m353 = m353 + 1) 
        begin: inbit353
            assign data_11[m353 + b353*16 + a12*28*16] = data_11_array[a12][b353][m353];
        end
    endgenerate
    generate 
        localparam integer b354 = 18;
        for (m354 = 0; m354 < 16; m354 = m354 + 1) 
        begin: inbit354
            assign data_11[m354 + b354*16 + a12*28*16] = data_11_array[a12][b354][m354];
        end
    endgenerate
    generate 
        localparam integer b355 = 19;
        for (m355 = 0; m355 < 16; m355 = m355 + 1) 
        begin: inbit355
            assign data_11[m355 + b355*16 + a12*28*16] = data_11_array[a12][b355][m355];
        end
    endgenerate
    generate 
        localparam integer b356 = 20;
        for (m356 = 0; m356 < 16; m356 = m356 + 1) 
        begin: inbit356
            assign data_11[m356 + b356*16 + a12*28*16] = data_11_array[a12][b356][m356];
        end
    endgenerate
    generate 
        localparam integer b357 = 21;
        for (m357 = 0; m357 < 16; m357 = m357 + 1) 
        begin: inbit357
            assign data_11[m357 + b357*16 + a12*28*16] = data_11_array[a12][b357][m357];
        end
    endgenerate
    generate 
        localparam integer b358 = 22;
        for (m358 = 0; m358 < 16; m358 = m358 + 1) 
        begin: inbit358
            assign data_11[m358 + b358*16 + a12*28*16] = data_11_array[a12][b358][m358];
        end
    endgenerate
    generate 
        localparam integer b359 = 23;
        for (m359 = 0; m359 < 16; m359 = m359 + 1) 
        begin: inbit359
            assign data_11[m359 + b359*16 + a12*28*16] = data_11_array[a12][b359][m359];
        end
    endgenerate
    generate 
        localparam integer b360 = 24;
        for (m360 = 0; m360 < 16; m360 = m360 + 1) 
        begin: inbit360
            assign data_11[m360 + b360*16 + a12*28*16] = data_11_array[a12][b360][m360];
        end
    endgenerate
    generate 
        localparam integer b361 = 25;
        for (m361 = 0; m361 < 16; m361 = m361 + 1) 
        begin: inbit361
            assign data_11[m361 + b361*16 + a12*28*16] = data_11_array[a12][b361][m361];
        end
    endgenerate
    generate 
        localparam integer b362 = 26;
        for (m362 = 0; m362 < 16; m362 = m362 + 1) 
        begin: inbit362
            assign data_11[m362 + b362*16 + a12*28*16] = data_11_array[a12][b362][m362];
        end
    endgenerate
    generate 
        localparam integer b363 = 27;
        for (m363 = 0; m363 < 16; m363 = m363 + 1) 
        begin: inbit363
            assign data_11[m363 + b363*16 + a12*28*16] = data_11_array[a12][b363][m363];
        end
    endgenerate
    localparam integer a13 = 13;
    generate 
        localparam integer b364 = 0;
        for (m364 = 0; m364 < 16; m364 = m364 + 1) 
        begin: inbit364
            assign data_11[m364 + b364*16 + a13*28*16] = data_11_array[a13][b364][m364];
        end
    endgenerate
    generate 
        localparam integer b365 = 1;
        for (m365 = 0; m365 < 16; m365 = m365 + 1) 
        begin: inbit365
            assign data_11[m365 + b365*16 + a13*28*16] = data_11_array[a13][b365][m365];
        end
    endgenerate
    generate 
        localparam integer b366 = 2;
        for (m366 = 0; m366 < 16; m366 = m366 + 1) 
        begin: inbit366
            assign data_11[m366 + b366*16 + a13*28*16] = data_11_array[a13][b366][m366];
        end
    endgenerate
    generate 
        localparam integer b367 = 3;
        for (m367 = 0; m367 < 16; m367 = m367 + 1) 
        begin: inbit367
            assign data_11[m367 + b367*16 + a13*28*16] = data_11_array[a13][b367][m367];
        end
    endgenerate
    generate 
        localparam integer b368 = 4;
        for (m368 = 0; m368 < 16; m368 = m368 + 1) 
        begin: inbit368
            assign data_11[m368 + b368*16 + a13*28*16] = data_11_array[a13][b368][m368];
        end
    endgenerate
    generate 
        localparam integer b369 = 5;
        for (m369 = 0; m369 < 16; m369 = m369 + 1) 
        begin: inbit369
            assign data_11[m369 + b369*16 + a13*28*16] = data_11_array[a13][b369][m369];
        end
    endgenerate
    generate 
        localparam integer b370 = 6;
        for (m370 = 0; m370 < 16; m370 = m370 + 1) 
        begin: inbit370
            assign data_11[m370 + b370*16 + a13*28*16] = data_11_array[a13][b370][m370];
        end
    endgenerate
    generate 
        localparam integer b371 = 7;
        for (m371 = 0; m371 < 16; m371 = m371 + 1) 
        begin: inbit371
            assign data_11[m371 + b371*16 + a13*28*16] = data_11_array[a13][b371][m371];
        end
    endgenerate
    generate 
        localparam integer b372 = 8;
        for (m372 = 0; m372 < 16; m372 = m372 + 1) 
        begin: inbit372
            assign data_11[m372 + b372*16 + a13*28*16] = data_11_array[a13][b372][m372];
        end
    endgenerate
    generate 
        localparam integer b373 = 9;
        for (m373 = 0; m373 < 16; m373 = m373 + 1) 
        begin: inbit373
            assign data_11[m373 + b373*16 + a13*28*16] = data_11_array[a13][b373][m373];
        end
    endgenerate
    generate 
        localparam integer b374 = 10;
        for (m374 = 0; m374 < 16; m374 = m374 + 1) 
        begin: inbit374
            assign data_11[m374 + b374*16 + a13*28*16] = data_11_array[a13][b374][m374];
        end
    endgenerate
    generate 
        localparam integer b375 = 11;
        for (m375 = 0; m375 < 16; m375 = m375 + 1) 
        begin: inbit375
            assign data_11[m375 + b375*16 + a13*28*16] = data_11_array[a13][b375][m375];
        end
    endgenerate
    generate 
        localparam integer b376 = 12;
        for (m376 = 0; m376 < 16; m376 = m376 + 1) 
        begin: inbit376
            assign data_11[m376 + b376*16 + a13*28*16] = data_11_array[a13][b376][m376];
        end
    endgenerate
    generate 
        localparam integer b377 = 13;
        for (m377 = 0; m377 < 16; m377 = m377 + 1) 
        begin: inbit377
            assign data_11[m377 + b377*16 + a13*28*16] = data_11_array[a13][b377][m377];
        end
    endgenerate
    generate 
        localparam integer b378 = 14;
        for (m378 = 0; m378 < 16; m378 = m378 + 1) 
        begin: inbit378
            assign data_11[m378 + b378*16 + a13*28*16] = data_11_array[a13][b378][m378];
        end
    endgenerate
    generate 
        localparam integer b379 = 15;
        for (m379 = 0; m379 < 16; m379 = m379 + 1) 
        begin: inbit379
            assign data_11[m379 + b379*16 + a13*28*16] = data_11_array[a13][b379][m379];
        end
    endgenerate
    generate 
        localparam integer b380 = 16;
        for (m380 = 0; m380 < 16; m380 = m380 + 1) 
        begin: inbit380
            assign data_11[m380 + b380*16 + a13*28*16] = data_11_array[a13][b380][m380];
        end
    endgenerate
    generate 
        localparam integer b381 = 17;
        for (m381 = 0; m381 < 16; m381 = m381 + 1) 
        begin: inbit381
            assign data_11[m381 + b381*16 + a13*28*16] = data_11_array[a13][b381][m381];
        end
    endgenerate
    generate 
        localparam integer b382 = 18;
        for (m382 = 0; m382 < 16; m382 = m382 + 1) 
        begin: inbit382
            assign data_11[m382 + b382*16 + a13*28*16] = data_11_array[a13][b382][m382];
        end
    endgenerate
    generate 
        localparam integer b383 = 19;
        for (m383 = 0; m383 < 16; m383 = m383 + 1) 
        begin: inbit383
            assign data_11[m383 + b383*16 + a13*28*16] = data_11_array[a13][b383][m383];
        end
    endgenerate
    generate 
        localparam integer b384 = 20;
        for (m384 = 0; m384 < 16; m384 = m384 + 1) 
        begin: inbit384
            assign data_11[m384 + b384*16 + a13*28*16] = data_11_array[a13][b384][m384];
        end
    endgenerate
    generate 
        localparam integer b385 = 21;
        for (m385 = 0; m385 < 16; m385 = m385 + 1) 
        begin: inbit385
            assign data_11[m385 + b385*16 + a13*28*16] = data_11_array[a13][b385][m385];
        end
    endgenerate
    generate 
        localparam integer b386 = 22;
        for (m386 = 0; m386 < 16; m386 = m386 + 1) 
        begin: inbit386
            assign data_11[m386 + b386*16 + a13*28*16] = data_11_array[a13][b386][m386];
        end
    endgenerate
    generate 
        localparam integer b387 = 23;
        for (m387 = 0; m387 < 16; m387 = m387 + 1) 
        begin: inbit387
            assign data_11[m387 + b387*16 + a13*28*16] = data_11_array[a13][b387][m387];
        end
    endgenerate
    generate 
        localparam integer b388 = 24;
        for (m388 = 0; m388 < 16; m388 = m388 + 1) 
        begin: inbit388
            assign data_11[m388 + b388*16 + a13*28*16] = data_11_array[a13][b388][m388];
        end
    endgenerate
    generate 
        localparam integer b389 = 25;
        for (m389 = 0; m389 < 16; m389 = m389 + 1) 
        begin: inbit389
            assign data_11[m389 + b389*16 + a13*28*16] = data_11_array[a13][b389][m389];
        end
    endgenerate
    generate 
        localparam integer b390 = 26;
        for (m390 = 0; m390 < 16; m390 = m390 + 1) 
        begin: inbit390
            assign data_11[m390 + b390*16 + a13*28*16] = data_11_array[a13][b390][m390];
        end
    endgenerate
    generate 
        localparam integer b391 = 27;
        for (m391 = 0; m391 < 16; m391 = m391 + 1) 
        begin: inbit391
            assign data_11[m391 + b391*16 + a13*28*16] = data_11_array[a13][b391][m391];
        end
    endgenerate
    localparam integer a14 = 14;
    generate 
        localparam integer b392 = 0;
        for (m392 = 0; m392 < 16; m392 = m392 + 1) 
        begin: inbit392
            assign data_11[m392 + b392*16 + a14*28*16] = data_11_array[a14][b392][m392];
        end
    endgenerate
    generate 
        localparam integer b393 = 1;
        for (m393 = 0; m393 < 16; m393 = m393 + 1) 
        begin: inbit393
            assign data_11[m393 + b393*16 + a14*28*16] = data_11_array[a14][b393][m393];
        end
    endgenerate
    generate 
        localparam integer b394 = 2;
        for (m394 = 0; m394 < 16; m394 = m394 + 1) 
        begin: inbit394
            assign data_11[m394 + b394*16 + a14*28*16] = data_11_array[a14][b394][m394];
        end
    endgenerate
    generate 
        localparam integer b395 = 3;
        for (m395 = 0; m395 < 16; m395 = m395 + 1) 
        begin: inbit395
            assign data_11[m395 + b395*16 + a14*28*16] = data_11_array[a14][b395][m395];
        end
    endgenerate
    generate 
        localparam integer b396 = 4;
        for (m396 = 0; m396 < 16; m396 = m396 + 1) 
        begin: inbit396
            assign data_11[m396 + b396*16 + a14*28*16] = data_11_array[a14][b396][m396];
        end
    endgenerate
    generate 
        localparam integer b397 = 5;
        for (m397 = 0; m397 < 16; m397 = m397 + 1) 
        begin: inbit397
            assign data_11[m397 + b397*16 + a14*28*16] = data_11_array[a14][b397][m397];
        end
    endgenerate
    generate 
        localparam integer b398 = 6;
        for (m398 = 0; m398 < 16; m398 = m398 + 1) 
        begin: inbit398
            assign data_11[m398 + b398*16 + a14*28*16] = data_11_array[a14][b398][m398];
        end
    endgenerate
    generate 
        localparam integer b399 = 7;
        for (m399 = 0; m399 < 16; m399 = m399 + 1) 
        begin: inbit399
            assign data_11[m399 + b399*16 + a14*28*16] = data_11_array[a14][b399][m399];
        end
    endgenerate
    generate 
        localparam integer b400 = 8;
        for (m400 = 0; m400 < 16; m400 = m400 + 1) 
        begin: inbit400
            assign data_11[m400 + b400*16 + a14*28*16] = data_11_array[a14][b400][m400];
        end
    endgenerate
    generate 
        localparam integer b401 = 9;
        for (m401 = 0; m401 < 16; m401 = m401 + 1) 
        begin: inbit401
            assign data_11[m401 + b401*16 + a14*28*16] = data_11_array[a14][b401][m401];
        end
    endgenerate
    generate 
        localparam integer b402 = 10;
        for (m402 = 0; m402 < 16; m402 = m402 + 1) 
        begin: inbit402
            assign data_11[m402 + b402*16 + a14*28*16] = data_11_array[a14][b402][m402];
        end
    endgenerate
    generate 
        localparam integer b403 = 11;
        for (m403 = 0; m403 < 16; m403 = m403 + 1) 
        begin: inbit403
            assign data_11[m403 + b403*16 + a14*28*16] = data_11_array[a14][b403][m403];
        end
    endgenerate
    generate 
        localparam integer b404 = 12;
        for (m404 = 0; m404 < 16; m404 = m404 + 1) 
        begin: inbit404
            assign data_11[m404 + b404*16 + a14*28*16] = data_11_array[a14][b404][m404];
        end
    endgenerate
    generate 
        localparam integer b405 = 13;
        for (m405 = 0; m405 < 16; m405 = m405 + 1) 
        begin: inbit405
            assign data_11[m405 + b405*16 + a14*28*16] = data_11_array[a14][b405][m405];
        end
    endgenerate
    generate 
        localparam integer b406 = 14;
        for (m406 = 0; m406 < 16; m406 = m406 + 1) 
        begin: inbit406
            assign data_11[m406 + b406*16 + a14*28*16] = data_11_array[a14][b406][m406];
        end
    endgenerate
    generate 
        localparam integer b407 = 15;
        for (m407 = 0; m407 < 16; m407 = m407 + 1) 
        begin: inbit407
            assign data_11[m407 + b407*16 + a14*28*16] = data_11_array[a14][b407][m407];
        end
    endgenerate
    generate 
        localparam integer b408 = 16;
        for (m408 = 0; m408 < 16; m408 = m408 + 1) 
        begin: inbit408
            assign data_11[m408 + b408*16 + a14*28*16] = data_11_array[a14][b408][m408];
        end
    endgenerate
    generate 
        localparam integer b409 = 17;
        for (m409 = 0; m409 < 16; m409 = m409 + 1) 
        begin: inbit409
            assign data_11[m409 + b409*16 + a14*28*16] = data_11_array[a14][b409][m409];
        end
    endgenerate
    generate 
        localparam integer b410 = 18;
        for (m410 = 0; m410 < 16; m410 = m410 + 1) 
        begin: inbit410
            assign data_11[m410 + b410*16 + a14*28*16] = data_11_array[a14][b410][m410];
        end
    endgenerate
    generate 
        localparam integer b411 = 19;
        for (m411 = 0; m411 < 16; m411 = m411 + 1) 
        begin: inbit411
            assign data_11[m411 + b411*16 + a14*28*16] = data_11_array[a14][b411][m411];
        end
    endgenerate
    generate 
        localparam integer b412 = 20;
        for (m412 = 0; m412 < 16; m412 = m412 + 1) 
        begin: inbit412
            assign data_11[m412 + b412*16 + a14*28*16] = data_11_array[a14][b412][m412];
        end
    endgenerate
    generate 
        localparam integer b413 = 21;
        for (m413 = 0; m413 < 16; m413 = m413 + 1) 
        begin: inbit413
            assign data_11[m413 + b413*16 + a14*28*16] = data_11_array[a14][b413][m413];
        end
    endgenerate
    generate 
        localparam integer b414 = 22;
        for (m414 = 0; m414 < 16; m414 = m414 + 1) 
        begin: inbit414
            assign data_11[m414 + b414*16 + a14*28*16] = data_11_array[a14][b414][m414];
        end
    endgenerate
    generate 
        localparam integer b415 = 23;
        for (m415 = 0; m415 < 16; m415 = m415 + 1) 
        begin: inbit415
            assign data_11[m415 + b415*16 + a14*28*16] = data_11_array[a14][b415][m415];
        end
    endgenerate
    generate 
        localparam integer b416 = 24;
        for (m416 = 0; m416 < 16; m416 = m416 + 1) 
        begin: inbit416
            assign data_11[m416 + b416*16 + a14*28*16] = data_11_array[a14][b416][m416];
        end
    endgenerate
    generate 
        localparam integer b417 = 25;
        for (m417 = 0; m417 < 16; m417 = m417 + 1) 
        begin: inbit417
            assign data_11[m417 + b417*16 + a14*28*16] = data_11_array[a14][b417][m417];
        end
    endgenerate
    generate 
        localparam integer b418 = 26;
        for (m418 = 0; m418 < 16; m418 = m418 + 1) 
        begin: inbit418
            assign data_11[m418 + b418*16 + a14*28*16] = data_11_array[a14][b418][m418];
        end
    endgenerate
    generate 
        localparam integer b419 = 27;
        for (m419 = 0; m419 < 16; m419 = m419 + 1) 
        begin: inbit419
            assign data_11[m419 + b419*16 + a14*28*16] = data_11_array[a14][b419][m419];
        end
    endgenerate
    localparam integer a15 = 15;
    generate 
        localparam integer b420 = 0;
        for (m420 = 0; m420 < 16; m420 = m420 + 1) 
        begin: inbit420
            assign data_11[m420 + b420*16 + a15*28*16] = data_11_array[a15][b420][m420];
        end
    endgenerate
    generate 
        localparam integer b421 = 1;
        for (m421 = 0; m421 < 16; m421 = m421 + 1) 
        begin: inbit421
            assign data_11[m421 + b421*16 + a15*28*16] = data_11_array[a15][b421][m421];
        end
    endgenerate
    generate 
        localparam integer b422 = 2;
        for (m422 = 0; m422 < 16; m422 = m422 + 1) 
        begin: inbit422
            assign data_11[m422 + b422*16 + a15*28*16] = data_11_array[a15][b422][m422];
        end
    endgenerate
    generate 
        localparam integer b423 = 3;
        for (m423 = 0; m423 < 16; m423 = m423 + 1) 
        begin: inbit423
            assign data_11[m423 + b423*16 + a15*28*16] = data_11_array[a15][b423][m423];
        end
    endgenerate
    generate 
        localparam integer b424 = 4;
        for (m424 = 0; m424 < 16; m424 = m424 + 1) 
        begin: inbit424
            assign data_11[m424 + b424*16 + a15*28*16] = data_11_array[a15][b424][m424];
        end
    endgenerate
    generate 
        localparam integer b425 = 5;
        for (m425 = 0; m425 < 16; m425 = m425 + 1) 
        begin: inbit425
            assign data_11[m425 + b425*16 + a15*28*16] = data_11_array[a15][b425][m425];
        end
    endgenerate
    generate 
        localparam integer b426 = 6;
        for (m426 = 0; m426 < 16; m426 = m426 + 1) 
        begin: inbit426
            assign data_11[m426 + b426*16 + a15*28*16] = data_11_array[a15][b426][m426];
        end
    endgenerate
    generate 
        localparam integer b427 = 7;
        for (m427 = 0; m427 < 16; m427 = m427 + 1) 
        begin: inbit427
            assign data_11[m427 + b427*16 + a15*28*16] = data_11_array[a15][b427][m427];
        end
    endgenerate
    generate 
        localparam integer b428 = 8;
        for (m428 = 0; m428 < 16; m428 = m428 + 1) 
        begin: inbit428
            assign data_11[m428 + b428*16 + a15*28*16] = data_11_array[a15][b428][m428];
        end
    endgenerate
    generate 
        localparam integer b429 = 9;
        for (m429 = 0; m429 < 16; m429 = m429 + 1) 
        begin: inbit429
            assign data_11[m429 + b429*16 + a15*28*16] = data_11_array[a15][b429][m429];
        end
    endgenerate
    generate 
        localparam integer b430 = 10;
        for (m430 = 0; m430 < 16; m430 = m430 + 1) 
        begin: inbit430
            assign data_11[m430 + b430*16 + a15*28*16] = data_11_array[a15][b430][m430];
        end
    endgenerate
    generate 
        localparam integer b431 = 11;
        for (m431 = 0; m431 < 16; m431 = m431 + 1) 
        begin: inbit431
            assign data_11[m431 + b431*16 + a15*28*16] = data_11_array[a15][b431][m431];
        end
    endgenerate
    generate 
        localparam integer b432 = 12;
        for (m432 = 0; m432 < 16; m432 = m432 + 1) 
        begin: inbit432
            assign data_11[m432 + b432*16 + a15*28*16] = data_11_array[a15][b432][m432];
        end
    endgenerate
    generate 
        localparam integer b433 = 13;
        for (m433 = 0; m433 < 16; m433 = m433 + 1) 
        begin: inbit433
            assign data_11[m433 + b433*16 + a15*28*16] = data_11_array[a15][b433][m433];
        end
    endgenerate
    generate 
        localparam integer b434 = 14;
        for (m434 = 0; m434 < 16; m434 = m434 + 1) 
        begin: inbit434
            assign data_11[m434 + b434*16 + a15*28*16] = data_11_array[a15][b434][m434];
        end
    endgenerate
    generate 
        localparam integer b435 = 15;
        for (m435 = 0; m435 < 16; m435 = m435 + 1) 
        begin: inbit435
            assign data_11[m435 + b435*16 + a15*28*16] = data_11_array[a15][b435][m435];
        end
    endgenerate
    generate 
        localparam integer b436 = 16;
        for (m436 = 0; m436 < 16; m436 = m436 + 1) 
        begin: inbit436
            assign data_11[m436 + b436*16 + a15*28*16] = data_11_array[a15][b436][m436];
        end
    endgenerate
    generate 
        localparam integer b437 = 17;
        for (m437 = 0; m437 < 16; m437 = m437 + 1) 
        begin: inbit437
            assign data_11[m437 + b437*16 + a15*28*16] = data_11_array[a15][b437][m437];
        end
    endgenerate
    generate 
        localparam integer b438 = 18;
        for (m438 = 0; m438 < 16; m438 = m438 + 1) 
        begin: inbit438
            assign data_11[m438 + b438*16 + a15*28*16] = data_11_array[a15][b438][m438];
        end
    endgenerate
    generate 
        localparam integer b439 = 19;
        for (m439 = 0; m439 < 16; m439 = m439 + 1) 
        begin: inbit439
            assign data_11[m439 + b439*16 + a15*28*16] = data_11_array[a15][b439][m439];
        end
    endgenerate
    generate 
        localparam integer b440 = 20;
        for (m440 = 0; m440 < 16; m440 = m440 + 1) 
        begin: inbit440
            assign data_11[m440 + b440*16 + a15*28*16] = data_11_array[a15][b440][m440];
        end
    endgenerate
    generate 
        localparam integer b441 = 21;
        for (m441 = 0; m441 < 16; m441 = m441 + 1) 
        begin: inbit441
            assign data_11[m441 + b441*16 + a15*28*16] = data_11_array[a15][b441][m441];
        end
    endgenerate
    generate 
        localparam integer b442 = 22;
        for (m442 = 0; m442 < 16; m442 = m442 + 1) 
        begin: inbit442
            assign data_11[m442 + b442*16 + a15*28*16] = data_11_array[a15][b442][m442];
        end
    endgenerate
    generate 
        localparam integer b443 = 23;
        for (m443 = 0; m443 < 16; m443 = m443 + 1) 
        begin: inbit443
            assign data_11[m443 + b443*16 + a15*28*16] = data_11_array[a15][b443][m443];
        end
    endgenerate
    generate 
        localparam integer b444 = 24;
        for (m444 = 0; m444 < 16; m444 = m444 + 1) 
        begin: inbit444
            assign data_11[m444 + b444*16 + a15*28*16] = data_11_array[a15][b444][m444];
        end
    endgenerate
    generate 
        localparam integer b445 = 25;
        for (m445 = 0; m445 < 16; m445 = m445 + 1) 
        begin: inbit445
            assign data_11[m445 + b445*16 + a15*28*16] = data_11_array[a15][b445][m445];
        end
    endgenerate
    generate 
        localparam integer b446 = 26;
        for (m446 = 0; m446 < 16; m446 = m446 + 1) 
        begin: inbit446
            assign data_11[m446 + b446*16 + a15*28*16] = data_11_array[a15][b446][m446];
        end
    endgenerate
    generate 
        localparam integer b447 = 27;
        for (m447 = 0; m447 < 16; m447 = m447 + 1) 
        begin: inbit447
            assign data_11[m447 + b447*16 + a15*28*16] = data_11_array[a15][b447][m447];
        end
    endgenerate
    localparam integer a16 = 16;
    generate 
        localparam integer b448 = 0;
        for (m448 = 0; m448 < 16; m448 = m448 + 1) 
        begin: inbit448
            assign data_11[m448 + b448*16 + a16*28*16] = data_11_array[a16][b448][m448];
        end
    endgenerate
    generate 
        localparam integer b449 = 1;
        for (m449 = 0; m449 < 16; m449 = m449 + 1) 
        begin: inbit449
            assign data_11[m449 + b449*16 + a16*28*16] = data_11_array[a16][b449][m449];
        end
    endgenerate
    generate 
        localparam integer b450 = 2;
        for (m450 = 0; m450 < 16; m450 = m450 + 1) 
        begin: inbit450
            assign data_11[m450 + b450*16 + a16*28*16] = data_11_array[a16][b450][m450];
        end
    endgenerate
    generate 
        localparam integer b451 = 3;
        for (m451 = 0; m451 < 16; m451 = m451 + 1) 
        begin: inbit451
            assign data_11[m451 + b451*16 + a16*28*16] = data_11_array[a16][b451][m451];
        end
    endgenerate
    generate 
        localparam integer b452 = 4;
        for (m452 = 0; m452 < 16; m452 = m452 + 1) 
        begin: inbit452
            assign data_11[m452 + b452*16 + a16*28*16] = data_11_array[a16][b452][m452];
        end
    endgenerate
    generate 
        localparam integer b453 = 5;
        for (m453 = 0; m453 < 16; m453 = m453 + 1) 
        begin: inbit453
            assign data_11[m453 + b453*16 + a16*28*16] = data_11_array[a16][b453][m453];
        end
    endgenerate
    generate 
        localparam integer b454 = 6;
        for (m454 = 0; m454 < 16; m454 = m454 + 1) 
        begin: inbit454
            assign data_11[m454 + b454*16 + a16*28*16] = data_11_array[a16][b454][m454];
        end
    endgenerate
    generate 
        localparam integer b455 = 7;
        for (m455 = 0; m455 < 16; m455 = m455 + 1) 
        begin: inbit455
            assign data_11[m455 + b455*16 + a16*28*16] = data_11_array[a16][b455][m455];
        end
    endgenerate
    generate 
        localparam integer b456 = 8;
        for (m456 = 0; m456 < 16; m456 = m456 + 1) 
        begin: inbit456
            assign data_11[m456 + b456*16 + a16*28*16] = data_11_array[a16][b456][m456];
        end
    endgenerate
    generate 
        localparam integer b457 = 9;
        for (m457 = 0; m457 < 16; m457 = m457 + 1) 
        begin: inbit457
            assign data_11[m457 + b457*16 + a16*28*16] = data_11_array[a16][b457][m457];
        end
    endgenerate
    generate 
        localparam integer b458 = 10;
        for (m458 = 0; m458 < 16; m458 = m458 + 1) 
        begin: inbit458
            assign data_11[m458 + b458*16 + a16*28*16] = data_11_array[a16][b458][m458];
        end
    endgenerate
    generate 
        localparam integer b459 = 11;
        for (m459 = 0; m459 < 16; m459 = m459 + 1) 
        begin: inbit459
            assign data_11[m459 + b459*16 + a16*28*16] = data_11_array[a16][b459][m459];
        end
    endgenerate
    generate 
        localparam integer b460 = 12;
        for (m460 = 0; m460 < 16; m460 = m460 + 1) 
        begin: inbit460
            assign data_11[m460 + b460*16 + a16*28*16] = data_11_array[a16][b460][m460];
        end
    endgenerate
    generate 
        localparam integer b461 = 13;
        for (m461 = 0; m461 < 16; m461 = m461 + 1) 
        begin: inbit461
            assign data_11[m461 + b461*16 + a16*28*16] = data_11_array[a16][b461][m461];
        end
    endgenerate
    generate 
        localparam integer b462 = 14;
        for (m462 = 0; m462 < 16; m462 = m462 + 1) 
        begin: inbit462
            assign data_11[m462 + b462*16 + a16*28*16] = data_11_array[a16][b462][m462];
        end
    endgenerate
    generate 
        localparam integer b463 = 15;
        for (m463 = 0; m463 < 16; m463 = m463 + 1) 
        begin: inbit463
            assign data_11[m463 + b463*16 + a16*28*16] = data_11_array[a16][b463][m463];
        end
    endgenerate
    generate 
        localparam integer b464 = 16;
        for (m464 = 0; m464 < 16; m464 = m464 + 1) 
        begin: inbit464
            assign data_11[m464 + b464*16 + a16*28*16] = data_11_array[a16][b464][m464];
        end
    endgenerate
    generate 
        localparam integer b465 = 17;
        for (m465 = 0; m465 < 16; m465 = m465 + 1) 
        begin: inbit465
            assign data_11[m465 + b465*16 + a16*28*16] = data_11_array[a16][b465][m465];
        end
    endgenerate
    generate 
        localparam integer b466 = 18;
        for (m466 = 0; m466 < 16; m466 = m466 + 1) 
        begin: inbit466
            assign data_11[m466 + b466*16 + a16*28*16] = data_11_array[a16][b466][m466];
        end
    endgenerate
    generate 
        localparam integer b467 = 19;
        for (m467 = 0; m467 < 16; m467 = m467 + 1) 
        begin: inbit467
            assign data_11[m467 + b467*16 + a16*28*16] = data_11_array[a16][b467][m467];
        end
    endgenerate
    generate 
        localparam integer b468 = 20;
        for (m468 = 0; m468 < 16; m468 = m468 + 1) 
        begin: inbit468
            assign data_11[m468 + b468*16 + a16*28*16] = data_11_array[a16][b468][m468];
        end
    endgenerate
    generate 
        localparam integer b469 = 21;
        for (m469 = 0; m469 < 16; m469 = m469 + 1) 
        begin: inbit469
            assign data_11[m469 + b469*16 + a16*28*16] = data_11_array[a16][b469][m469];
        end
    endgenerate
    generate 
        localparam integer b470 = 22;
        for (m470 = 0; m470 < 16; m470 = m470 + 1) 
        begin: inbit470
            assign data_11[m470 + b470*16 + a16*28*16] = data_11_array[a16][b470][m470];
        end
    endgenerate
    generate 
        localparam integer b471 = 23;
        for (m471 = 0; m471 < 16; m471 = m471 + 1) 
        begin: inbit471
            assign data_11[m471 + b471*16 + a16*28*16] = data_11_array[a16][b471][m471];
        end
    endgenerate
    generate 
        localparam integer b472 = 24;
        for (m472 = 0; m472 < 16; m472 = m472 + 1) 
        begin: inbit472
            assign data_11[m472 + b472*16 + a16*28*16] = data_11_array[a16][b472][m472];
        end
    endgenerate
    generate 
        localparam integer b473 = 25;
        for (m473 = 0; m473 < 16; m473 = m473 + 1) 
        begin: inbit473
            assign data_11[m473 + b473*16 + a16*28*16] = data_11_array[a16][b473][m473];
        end
    endgenerate
    generate 
        localparam integer b474 = 26;
        for (m474 = 0; m474 < 16; m474 = m474 + 1) 
        begin: inbit474
            assign data_11[m474 + b474*16 + a16*28*16] = data_11_array[a16][b474][m474];
        end
    endgenerate
    generate 
        localparam integer b475 = 27;
        for (m475 = 0; m475 < 16; m475 = m475 + 1) 
        begin: inbit475
            assign data_11[m475 + b475*16 + a16*28*16] = data_11_array[a16][b475][m475];
        end
    endgenerate
    localparam integer a17 = 17;
    generate 
        localparam integer b476 = 0;
        for (m476 = 0; m476 < 16; m476 = m476 + 1) 
        begin: inbit476
            assign data_11[m476 + b476*16 + a17*28*16] = data_11_array[a17][b476][m476];
        end
    endgenerate
    generate 
        localparam integer b477 = 1;
        for (m477 = 0; m477 < 16; m477 = m477 + 1) 
        begin: inbit477
            assign data_11[m477 + b477*16 + a17*28*16] = data_11_array[a17][b477][m477];
        end
    endgenerate
    generate 
        localparam integer b478 = 2;
        for (m478 = 0; m478 < 16; m478 = m478 + 1) 
        begin: inbit478
            assign data_11[m478 + b478*16 + a17*28*16] = data_11_array[a17][b478][m478];
        end
    endgenerate
    generate 
        localparam integer b479 = 3;
        for (m479 = 0; m479 < 16; m479 = m479 + 1) 
        begin: inbit479
            assign data_11[m479 + b479*16 + a17*28*16] = data_11_array[a17][b479][m479];
        end
    endgenerate
    generate 
        localparam integer b480 = 4;
        for (m480 = 0; m480 < 16; m480 = m480 + 1) 
        begin: inbit480
            assign data_11[m480 + b480*16 + a17*28*16] = data_11_array[a17][b480][m480];
        end
    endgenerate
    generate 
        localparam integer b481 = 5;
        for (m481 = 0; m481 < 16; m481 = m481 + 1) 
        begin: inbit481
            assign data_11[m481 + b481*16 + a17*28*16] = data_11_array[a17][b481][m481];
        end
    endgenerate
    generate 
        localparam integer b482 = 6;
        for (m482 = 0; m482 < 16; m482 = m482 + 1) 
        begin: inbit482
            assign data_11[m482 + b482*16 + a17*28*16] = data_11_array[a17][b482][m482];
        end
    endgenerate
    generate 
        localparam integer b483 = 7;
        for (m483 = 0; m483 < 16; m483 = m483 + 1) 
        begin: inbit483
            assign data_11[m483 + b483*16 + a17*28*16] = data_11_array[a17][b483][m483];
        end
    endgenerate
    generate 
        localparam integer b484 = 8;
        for (m484 = 0; m484 < 16; m484 = m484 + 1) 
        begin: inbit484
            assign data_11[m484 + b484*16 + a17*28*16] = data_11_array[a17][b484][m484];
        end
    endgenerate
    generate 
        localparam integer b485 = 9;
        for (m485 = 0; m485 < 16; m485 = m485 + 1) 
        begin: inbit485
            assign data_11[m485 + b485*16 + a17*28*16] = data_11_array[a17][b485][m485];
        end
    endgenerate
    generate 
        localparam integer b486 = 10;
        for (m486 = 0; m486 < 16; m486 = m486 + 1) 
        begin: inbit486
            assign data_11[m486 + b486*16 + a17*28*16] = data_11_array[a17][b486][m486];
        end
    endgenerate
    generate 
        localparam integer b487 = 11;
        for (m487 = 0; m487 < 16; m487 = m487 + 1) 
        begin: inbit487
            assign data_11[m487 + b487*16 + a17*28*16] = data_11_array[a17][b487][m487];
        end
    endgenerate
    generate 
        localparam integer b488 = 12;
        for (m488 = 0; m488 < 16; m488 = m488 + 1) 
        begin: inbit488
            assign data_11[m488 + b488*16 + a17*28*16] = data_11_array[a17][b488][m488];
        end
    endgenerate
    generate 
        localparam integer b489 = 13;
        for (m489 = 0; m489 < 16; m489 = m489 + 1) 
        begin: inbit489
            assign data_11[m489 + b489*16 + a17*28*16] = data_11_array[a17][b489][m489];
        end
    endgenerate
    generate 
        localparam integer b490 = 14;
        for (m490 = 0; m490 < 16; m490 = m490 + 1) 
        begin: inbit490
            assign data_11[m490 + b490*16 + a17*28*16] = data_11_array[a17][b490][m490];
        end
    endgenerate
    generate 
        localparam integer b491 = 15;
        for (m491 = 0; m491 < 16; m491 = m491 + 1) 
        begin: inbit491
            assign data_11[m491 + b491*16 + a17*28*16] = data_11_array[a17][b491][m491];
        end
    endgenerate
    generate 
        localparam integer b492 = 16;
        for (m492 = 0; m492 < 16; m492 = m492 + 1) 
        begin: inbit492
            assign data_11[m492 + b492*16 + a17*28*16] = data_11_array[a17][b492][m492];
        end
    endgenerate
    generate 
        localparam integer b493 = 17;
        for (m493 = 0; m493 < 16; m493 = m493 + 1) 
        begin: inbit493
            assign data_11[m493 + b493*16 + a17*28*16] = data_11_array[a17][b493][m493];
        end
    endgenerate
    generate 
        localparam integer b494 = 18;
        for (m494 = 0; m494 < 16; m494 = m494 + 1) 
        begin: inbit494
            assign data_11[m494 + b494*16 + a17*28*16] = data_11_array[a17][b494][m494];
        end
    endgenerate
    generate 
        localparam integer b495 = 19;
        for (m495 = 0; m495 < 16; m495 = m495 + 1) 
        begin: inbit495
            assign data_11[m495 + b495*16 + a17*28*16] = data_11_array[a17][b495][m495];
        end
    endgenerate
    generate 
        localparam integer b496 = 20;
        for (m496 = 0; m496 < 16; m496 = m496 + 1) 
        begin: inbit496
            assign data_11[m496 + b496*16 + a17*28*16] = data_11_array[a17][b496][m496];
        end
    endgenerate
    generate 
        localparam integer b497 = 21;
        for (m497 = 0; m497 < 16; m497 = m497 + 1) 
        begin: inbit497
            assign data_11[m497 + b497*16 + a17*28*16] = data_11_array[a17][b497][m497];
        end
    endgenerate
    generate 
        localparam integer b498 = 22;
        for (m498 = 0; m498 < 16; m498 = m498 + 1) 
        begin: inbit498
            assign data_11[m498 + b498*16 + a17*28*16] = data_11_array[a17][b498][m498];
        end
    endgenerate
    generate 
        localparam integer b499 = 23;
        for (m499 = 0; m499 < 16; m499 = m499 + 1) 
        begin: inbit499
            assign data_11[m499 + b499*16 + a17*28*16] = data_11_array[a17][b499][m499];
        end
    endgenerate
    generate 
        localparam integer b500 = 24;
        for (m500 = 0; m500 < 16; m500 = m500 + 1) 
        begin: inbit500
            assign data_11[m500 + b500*16 + a17*28*16] = data_11_array[a17][b500][m500];
        end
    endgenerate
    generate 
        localparam integer b501 = 25;
        for (m501 = 0; m501 < 16; m501 = m501 + 1) 
        begin: inbit501
            assign data_11[m501 + b501*16 + a17*28*16] = data_11_array[a17][b501][m501];
        end
    endgenerate
    generate 
        localparam integer b502 = 26;
        for (m502 = 0; m502 < 16; m502 = m502 + 1) 
        begin: inbit502
            assign data_11[m502 + b502*16 + a17*28*16] = data_11_array[a17][b502][m502];
        end
    endgenerate
    generate 
        localparam integer b503 = 27;
        for (m503 = 0; m503 < 16; m503 = m503 + 1) 
        begin: inbit503
            assign data_11[m503 + b503*16 + a17*28*16] = data_11_array[a17][b503][m503];
        end
    endgenerate
    localparam integer a18 = 18;
    generate 
        localparam integer b504 = 0;
        for (m504 = 0; m504 < 16; m504 = m504 + 1) 
        begin: inbit504
            assign data_11[m504 + b504*16 + a18*28*16] = data_11_array[a18][b504][m504];
        end
    endgenerate
    generate 
        localparam integer b505 = 1;
        for (m505 = 0; m505 < 16; m505 = m505 + 1) 
        begin: inbit505
            assign data_11[m505 + b505*16 + a18*28*16] = data_11_array[a18][b505][m505];
        end
    endgenerate
    generate 
        localparam integer b506 = 2;
        for (m506 = 0; m506 < 16; m506 = m506 + 1) 
        begin: inbit506
            assign data_11[m506 + b506*16 + a18*28*16] = data_11_array[a18][b506][m506];
        end
    endgenerate
    generate 
        localparam integer b507 = 3;
        for (m507 = 0; m507 < 16; m507 = m507 + 1) 
        begin: inbit507
            assign data_11[m507 + b507*16 + a18*28*16] = data_11_array[a18][b507][m507];
        end
    endgenerate
    generate 
        localparam integer b508 = 4;
        for (m508 = 0; m508 < 16; m508 = m508 + 1) 
        begin: inbit508
            assign data_11[m508 + b508*16 + a18*28*16] = data_11_array[a18][b508][m508];
        end
    endgenerate
    generate 
        localparam integer b509 = 5;
        for (m509 = 0; m509 < 16; m509 = m509 + 1) 
        begin: inbit509
            assign data_11[m509 + b509*16 + a18*28*16] = data_11_array[a18][b509][m509];
        end
    endgenerate
    generate 
        localparam integer b510 = 6;
        for (m510 = 0; m510 < 16; m510 = m510 + 1) 
        begin: inbit510
            assign data_11[m510 + b510*16 + a18*28*16] = data_11_array[a18][b510][m510];
        end
    endgenerate
    generate 
        localparam integer b511 = 7;
        for (m511 = 0; m511 < 16; m511 = m511 + 1) 
        begin: inbit511
            assign data_11[m511 + b511*16 + a18*28*16] = data_11_array[a18][b511][m511];
        end
    endgenerate
    generate 
        localparam integer b512 = 8;
        for (m512 = 0; m512 < 16; m512 = m512 + 1) 
        begin: inbit512
            assign data_11[m512 + b512*16 + a18*28*16] = data_11_array[a18][b512][m512];
        end
    endgenerate
    generate 
        localparam integer b513 = 9;
        for (m513 = 0; m513 < 16; m513 = m513 + 1) 
        begin: inbit513
            assign data_11[m513 + b513*16 + a18*28*16] = data_11_array[a18][b513][m513];
        end
    endgenerate
    generate 
        localparam integer b514 = 10;
        for (m514 = 0; m514 < 16; m514 = m514 + 1) 
        begin: inbit514
            assign data_11[m514 + b514*16 + a18*28*16] = data_11_array[a18][b514][m514];
        end
    endgenerate
    generate 
        localparam integer b515 = 11;
        for (m515 = 0; m515 < 16; m515 = m515 + 1) 
        begin: inbit515
            assign data_11[m515 + b515*16 + a18*28*16] = data_11_array[a18][b515][m515];
        end
    endgenerate
    generate 
        localparam integer b516 = 12;
        for (m516 = 0; m516 < 16; m516 = m516 + 1) 
        begin: inbit516
            assign data_11[m516 + b516*16 + a18*28*16] = data_11_array[a18][b516][m516];
        end
    endgenerate
    generate 
        localparam integer b517 = 13;
        for (m517 = 0; m517 < 16; m517 = m517 + 1) 
        begin: inbit517
            assign data_11[m517 + b517*16 + a18*28*16] = data_11_array[a18][b517][m517];
        end
    endgenerate
    generate 
        localparam integer b518 = 14;
        for (m518 = 0; m518 < 16; m518 = m518 + 1) 
        begin: inbit518
            assign data_11[m518 + b518*16 + a18*28*16] = data_11_array[a18][b518][m518];
        end
    endgenerate
    generate 
        localparam integer b519 = 15;
        for (m519 = 0; m519 < 16; m519 = m519 + 1) 
        begin: inbit519
            assign data_11[m519 + b519*16 + a18*28*16] = data_11_array[a18][b519][m519];
        end
    endgenerate
    generate 
        localparam integer b520 = 16;
        for (m520 = 0; m520 < 16; m520 = m520 + 1) 
        begin: inbit520
            assign data_11[m520 + b520*16 + a18*28*16] = data_11_array[a18][b520][m520];
        end
    endgenerate
    generate 
        localparam integer b521 = 17;
        for (m521 = 0; m521 < 16; m521 = m521 + 1) 
        begin: inbit521
            assign data_11[m521 + b521*16 + a18*28*16] = data_11_array[a18][b521][m521];
        end
    endgenerate
    generate 
        localparam integer b522 = 18;
        for (m522 = 0; m522 < 16; m522 = m522 + 1) 
        begin: inbit522
            assign data_11[m522 + b522*16 + a18*28*16] = data_11_array[a18][b522][m522];
        end
    endgenerate
    generate 
        localparam integer b523 = 19;
        for (m523 = 0; m523 < 16; m523 = m523 + 1) 
        begin: inbit523
            assign data_11[m523 + b523*16 + a18*28*16] = data_11_array[a18][b523][m523];
        end
    endgenerate
    generate 
        localparam integer b524 = 20;
        for (m524 = 0; m524 < 16; m524 = m524 + 1) 
        begin: inbit524
            assign data_11[m524 + b524*16 + a18*28*16] = data_11_array[a18][b524][m524];
        end
    endgenerate
    generate 
        localparam integer b525 = 21;
        for (m525 = 0; m525 < 16; m525 = m525 + 1) 
        begin: inbit525
            assign data_11[m525 + b525*16 + a18*28*16] = data_11_array[a18][b525][m525];
        end
    endgenerate
    generate 
        localparam integer b526 = 22;
        for (m526 = 0; m526 < 16; m526 = m526 + 1) 
        begin: inbit526
            assign data_11[m526 + b526*16 + a18*28*16] = data_11_array[a18][b526][m526];
        end
    endgenerate
    generate 
        localparam integer b527 = 23;
        for (m527 = 0; m527 < 16; m527 = m527 + 1) 
        begin: inbit527
            assign data_11[m527 + b527*16 + a18*28*16] = data_11_array[a18][b527][m527];
        end
    endgenerate
    generate 
        localparam integer b528 = 24;
        for (m528 = 0; m528 < 16; m528 = m528 + 1) 
        begin: inbit528
            assign data_11[m528 + b528*16 + a18*28*16] = data_11_array[a18][b528][m528];
        end
    endgenerate
    generate 
        localparam integer b529 = 25;
        for (m529 = 0; m529 < 16; m529 = m529 + 1) 
        begin: inbit529
            assign data_11[m529 + b529*16 + a18*28*16] = data_11_array[a18][b529][m529];
        end
    endgenerate
    generate 
        localparam integer b530 = 26;
        for (m530 = 0; m530 < 16; m530 = m530 + 1) 
        begin: inbit530
            assign data_11[m530 + b530*16 + a18*28*16] = data_11_array[a18][b530][m530];
        end
    endgenerate
    generate 
        localparam integer b531 = 27;
        for (m531 = 0; m531 < 16; m531 = m531 + 1) 
        begin: inbit531
            assign data_11[m531 + b531*16 + a18*28*16] = data_11_array[a18][b531][m531];
        end
    endgenerate
    localparam integer a19 = 19;
    generate 
        localparam integer b532 = 0;
        for (m532 = 0; m532 < 16; m532 = m532 + 1) 
        begin: inbit532
            assign data_11[m532 + b532*16 + a19*28*16] = data_11_array[a19][b532][m532];
        end
    endgenerate
    generate 
        localparam integer b533 = 1;
        for (m533 = 0; m533 < 16; m533 = m533 + 1) 
        begin: inbit533
            assign data_11[m533 + b533*16 + a19*28*16] = data_11_array[a19][b533][m533];
        end
    endgenerate
    generate 
        localparam integer b534 = 2;
        for (m534 = 0; m534 < 16; m534 = m534 + 1) 
        begin: inbit534
            assign data_11[m534 + b534*16 + a19*28*16] = data_11_array[a19][b534][m534];
        end
    endgenerate
    generate 
        localparam integer b535 = 3;
        for (m535 = 0; m535 < 16; m535 = m535 + 1) 
        begin: inbit535
            assign data_11[m535 + b535*16 + a19*28*16] = data_11_array[a19][b535][m535];
        end
    endgenerate
    generate 
        localparam integer b536 = 4;
        for (m536 = 0; m536 < 16; m536 = m536 + 1) 
        begin: inbit536
            assign data_11[m536 + b536*16 + a19*28*16] = data_11_array[a19][b536][m536];
        end
    endgenerate
    generate 
        localparam integer b537 = 5;
        for (m537 = 0; m537 < 16; m537 = m537 + 1) 
        begin: inbit537
            assign data_11[m537 + b537*16 + a19*28*16] = data_11_array[a19][b537][m537];
        end
    endgenerate
    generate 
        localparam integer b538 = 6;
        for (m538 = 0; m538 < 16; m538 = m538 + 1) 
        begin: inbit538
            assign data_11[m538 + b538*16 + a19*28*16] = data_11_array[a19][b538][m538];
        end
    endgenerate
    generate 
        localparam integer b539 = 7;
        for (m539 = 0; m539 < 16; m539 = m539 + 1) 
        begin: inbit539
            assign data_11[m539 + b539*16 + a19*28*16] = data_11_array[a19][b539][m539];
        end
    endgenerate
    generate 
        localparam integer b540 = 8;
        for (m540 = 0; m540 < 16; m540 = m540 + 1) 
        begin: inbit540
            assign data_11[m540 + b540*16 + a19*28*16] = data_11_array[a19][b540][m540];
        end
    endgenerate
    generate 
        localparam integer b541 = 9;
        for (m541 = 0; m541 < 16; m541 = m541 + 1) 
        begin: inbit541
            assign data_11[m541 + b541*16 + a19*28*16] = data_11_array[a19][b541][m541];
        end
    endgenerate
    generate 
        localparam integer b542 = 10;
        for (m542 = 0; m542 < 16; m542 = m542 + 1) 
        begin: inbit542
            assign data_11[m542 + b542*16 + a19*28*16] = data_11_array[a19][b542][m542];
        end
    endgenerate
    generate 
        localparam integer b543 = 11;
        for (m543 = 0; m543 < 16; m543 = m543 + 1) 
        begin: inbit543
            assign data_11[m543 + b543*16 + a19*28*16] = data_11_array[a19][b543][m543];
        end
    endgenerate
    generate 
        localparam integer b544 = 12;
        for (m544 = 0; m544 < 16; m544 = m544 + 1) 
        begin: inbit544
            assign data_11[m544 + b544*16 + a19*28*16] = data_11_array[a19][b544][m544];
        end
    endgenerate
    generate 
        localparam integer b545 = 13;
        for (m545 = 0; m545 < 16; m545 = m545 + 1) 
        begin: inbit545
            assign data_11[m545 + b545*16 + a19*28*16] = data_11_array[a19][b545][m545];
        end
    endgenerate
    generate 
        localparam integer b546 = 14;
        for (m546 = 0; m546 < 16; m546 = m546 + 1) 
        begin: inbit546
            assign data_11[m546 + b546*16 + a19*28*16] = data_11_array[a19][b546][m546];
        end
    endgenerate
    generate 
        localparam integer b547 = 15;
        for (m547 = 0; m547 < 16; m547 = m547 + 1) 
        begin: inbit547
            assign data_11[m547 + b547*16 + a19*28*16] = data_11_array[a19][b547][m547];
        end
    endgenerate
    generate 
        localparam integer b548 = 16;
        for (m548 = 0; m548 < 16; m548 = m548 + 1) 
        begin: inbit548
            assign data_11[m548 + b548*16 + a19*28*16] = data_11_array[a19][b548][m548];
        end
    endgenerate
    generate 
        localparam integer b549 = 17;
        for (m549 = 0; m549 < 16; m549 = m549 + 1) 
        begin: inbit549
            assign data_11[m549 + b549*16 + a19*28*16] = data_11_array[a19][b549][m549];
        end
    endgenerate
    generate 
        localparam integer b550 = 18;
        for (m550 = 0; m550 < 16; m550 = m550 + 1) 
        begin: inbit550
            assign data_11[m550 + b550*16 + a19*28*16] = data_11_array[a19][b550][m550];
        end
    endgenerate
    generate 
        localparam integer b551 = 19;
        for (m551 = 0; m551 < 16; m551 = m551 + 1) 
        begin: inbit551
            assign data_11[m551 + b551*16 + a19*28*16] = data_11_array[a19][b551][m551];
        end
    endgenerate
    generate 
        localparam integer b552 = 20;
        for (m552 = 0; m552 < 16; m552 = m552 + 1) 
        begin: inbit552
            assign data_11[m552 + b552*16 + a19*28*16] = data_11_array[a19][b552][m552];
        end
    endgenerate
    generate 
        localparam integer b553 = 21;
        for (m553 = 0; m553 < 16; m553 = m553 + 1) 
        begin: inbit553
            assign data_11[m553 + b553*16 + a19*28*16] = data_11_array[a19][b553][m553];
        end
    endgenerate
    generate 
        localparam integer b554 = 22;
        for (m554 = 0; m554 < 16; m554 = m554 + 1) 
        begin: inbit554
            assign data_11[m554 + b554*16 + a19*28*16] = data_11_array[a19][b554][m554];
        end
    endgenerate
    generate 
        localparam integer b555 = 23;
        for (m555 = 0; m555 < 16; m555 = m555 + 1) 
        begin: inbit555
            assign data_11[m555 + b555*16 + a19*28*16] = data_11_array[a19][b555][m555];
        end
    endgenerate
    generate 
        localparam integer b556 = 24;
        for (m556 = 0; m556 < 16; m556 = m556 + 1) 
        begin: inbit556
            assign data_11[m556 + b556*16 + a19*28*16] = data_11_array[a19][b556][m556];
        end
    endgenerate
    generate 
        localparam integer b557 = 25;
        for (m557 = 0; m557 < 16; m557 = m557 + 1) 
        begin: inbit557
            assign data_11[m557 + b557*16 + a19*28*16] = data_11_array[a19][b557][m557];
        end
    endgenerate
    generate 
        localparam integer b558 = 26;
        for (m558 = 0; m558 < 16; m558 = m558 + 1) 
        begin: inbit558
            assign data_11[m558 + b558*16 + a19*28*16] = data_11_array[a19][b558][m558];
        end
    endgenerate
    generate 
        localparam integer b559 = 27;
        for (m559 = 0; m559 < 16; m559 = m559 + 1) 
        begin: inbit559
            assign data_11[m559 + b559*16 + a19*28*16] = data_11_array[a19][b559][m559];
        end
    endgenerate
    localparam integer a20 = 20;
    generate 
        localparam integer b560 = 0;
        for (m560 = 0; m560 < 16; m560 = m560 + 1) 
        begin: inbit560
            assign data_11[m560 + b560*16 + a20*28*16] = data_11_array[a20][b560][m560];
        end
    endgenerate
    generate 
        localparam integer b561 = 1;
        for (m561 = 0; m561 < 16; m561 = m561 + 1) 
        begin: inbit561
            assign data_11[m561 + b561*16 + a20*28*16] = data_11_array[a20][b561][m561];
        end
    endgenerate
    generate 
        localparam integer b562 = 2;
        for (m562 = 0; m562 < 16; m562 = m562 + 1) 
        begin: inbit562
            assign data_11[m562 + b562*16 + a20*28*16] = data_11_array[a20][b562][m562];
        end
    endgenerate
    generate 
        localparam integer b563 = 3;
        for (m563 = 0; m563 < 16; m563 = m563 + 1) 
        begin: inbit563
            assign data_11[m563 + b563*16 + a20*28*16] = data_11_array[a20][b563][m563];
        end
    endgenerate
    generate 
        localparam integer b564 = 4;
        for (m564 = 0; m564 < 16; m564 = m564 + 1) 
        begin: inbit564
            assign data_11[m564 + b564*16 + a20*28*16] = data_11_array[a20][b564][m564];
        end
    endgenerate
    generate 
        localparam integer b565 = 5;
        for (m565 = 0; m565 < 16; m565 = m565 + 1) 
        begin: inbit565
            assign data_11[m565 + b565*16 + a20*28*16] = data_11_array[a20][b565][m565];
        end
    endgenerate
    generate 
        localparam integer b566 = 6;
        for (m566 = 0; m566 < 16; m566 = m566 + 1) 
        begin: inbit566
            assign data_11[m566 + b566*16 + a20*28*16] = data_11_array[a20][b566][m566];
        end
    endgenerate
    generate 
        localparam integer b567 = 7;
        for (m567 = 0; m567 < 16; m567 = m567 + 1) 
        begin: inbit567
            assign data_11[m567 + b567*16 + a20*28*16] = data_11_array[a20][b567][m567];
        end
    endgenerate
    generate 
        localparam integer b568 = 8;
        for (m568 = 0; m568 < 16; m568 = m568 + 1) 
        begin: inbit568
            assign data_11[m568 + b568*16 + a20*28*16] = data_11_array[a20][b568][m568];
        end
    endgenerate
    generate 
        localparam integer b569 = 9;
        for (m569 = 0; m569 < 16; m569 = m569 + 1) 
        begin: inbit569
            assign data_11[m569 + b569*16 + a20*28*16] = data_11_array[a20][b569][m569];
        end
    endgenerate
    generate 
        localparam integer b570 = 10;
        for (m570 = 0; m570 < 16; m570 = m570 + 1) 
        begin: inbit570
            assign data_11[m570 + b570*16 + a20*28*16] = data_11_array[a20][b570][m570];
        end
    endgenerate
    generate 
        localparam integer b571 = 11;
        for (m571 = 0; m571 < 16; m571 = m571 + 1) 
        begin: inbit571
            assign data_11[m571 + b571*16 + a20*28*16] = data_11_array[a20][b571][m571];
        end
    endgenerate
    generate 
        localparam integer b572 = 12;
        for (m572 = 0; m572 < 16; m572 = m572 + 1) 
        begin: inbit572
            assign data_11[m572 + b572*16 + a20*28*16] = data_11_array[a20][b572][m572];
        end
    endgenerate
    generate 
        localparam integer b573 = 13;
        for (m573 = 0; m573 < 16; m573 = m573 + 1) 
        begin: inbit573
            assign data_11[m573 + b573*16 + a20*28*16] = data_11_array[a20][b573][m573];
        end
    endgenerate
    generate 
        localparam integer b574 = 14;
        for (m574 = 0; m574 < 16; m574 = m574 + 1) 
        begin: inbit574
            assign data_11[m574 + b574*16 + a20*28*16] = data_11_array[a20][b574][m574];
        end
    endgenerate
    generate 
        localparam integer b575 = 15;
        for (m575 = 0; m575 < 16; m575 = m575 + 1) 
        begin: inbit575
            assign data_11[m575 + b575*16 + a20*28*16] = data_11_array[a20][b575][m575];
        end
    endgenerate
    generate 
        localparam integer b576 = 16;
        for (m576 = 0; m576 < 16; m576 = m576 + 1) 
        begin: inbit576
            assign data_11[m576 + b576*16 + a20*28*16] = data_11_array[a20][b576][m576];
        end
    endgenerate
    generate 
        localparam integer b577 = 17;
        for (m577 = 0; m577 < 16; m577 = m577 + 1) 
        begin: inbit577
            assign data_11[m577 + b577*16 + a20*28*16] = data_11_array[a20][b577][m577];
        end
    endgenerate
    generate 
        localparam integer b578 = 18;
        for (m578 = 0; m578 < 16; m578 = m578 + 1) 
        begin: inbit578
            assign data_11[m578 + b578*16 + a20*28*16] = data_11_array[a20][b578][m578];
        end
    endgenerate
    generate 
        localparam integer b579 = 19;
        for (m579 = 0; m579 < 16; m579 = m579 + 1) 
        begin: inbit579
            assign data_11[m579 + b579*16 + a20*28*16] = data_11_array[a20][b579][m579];
        end
    endgenerate
    generate 
        localparam integer b580 = 20;
        for (m580 = 0; m580 < 16; m580 = m580 + 1) 
        begin: inbit580
            assign data_11[m580 + b580*16 + a20*28*16] = data_11_array[a20][b580][m580];
        end
    endgenerate
    generate 
        localparam integer b581 = 21;
        for (m581 = 0; m581 < 16; m581 = m581 + 1) 
        begin: inbit581
            assign data_11[m581 + b581*16 + a20*28*16] = data_11_array[a20][b581][m581];
        end
    endgenerate
    generate 
        localparam integer b582 = 22;
        for (m582 = 0; m582 < 16; m582 = m582 + 1) 
        begin: inbit582
            assign data_11[m582 + b582*16 + a20*28*16] = data_11_array[a20][b582][m582];
        end
    endgenerate
    generate 
        localparam integer b583 = 23;
        for (m583 = 0; m583 < 16; m583 = m583 + 1) 
        begin: inbit583
            assign data_11[m583 + b583*16 + a20*28*16] = data_11_array[a20][b583][m583];
        end
    endgenerate
    generate 
        localparam integer b584 = 24;
        for (m584 = 0; m584 < 16; m584 = m584 + 1) 
        begin: inbit584
            assign data_11[m584 + b584*16 + a20*28*16] = data_11_array[a20][b584][m584];
        end
    endgenerate
    generate 
        localparam integer b585 = 25;
        for (m585 = 0; m585 < 16; m585 = m585 + 1) 
        begin: inbit585
            assign data_11[m585 + b585*16 + a20*28*16] = data_11_array[a20][b585][m585];
        end
    endgenerate
    generate 
        localparam integer b586 = 26;
        for (m586 = 0; m586 < 16; m586 = m586 + 1) 
        begin: inbit586
            assign data_11[m586 + b586*16 + a20*28*16] = data_11_array[a20][b586][m586];
        end
    endgenerate
    generate 
        localparam integer b587 = 27;
        for (m587 = 0; m587 < 16; m587 = m587 + 1) 
        begin: inbit587
            assign data_11[m587 + b587*16 + a20*28*16] = data_11_array[a20][b587][m587];
        end
    endgenerate
    localparam integer a21 = 21;
    generate 
        localparam integer b588 = 0;
        for (m588 = 0; m588 < 16; m588 = m588 + 1) 
        begin: inbit588
            assign data_11[m588 + b588*16 + a21*28*16] = data_11_array[a21][b588][m588];
        end
    endgenerate
    generate 
        localparam integer b589 = 1;
        for (m589 = 0; m589 < 16; m589 = m589 + 1) 
        begin: inbit589
            assign data_11[m589 + b589*16 + a21*28*16] = data_11_array[a21][b589][m589];
        end
    endgenerate
    generate 
        localparam integer b590 = 2;
        for (m590 = 0; m590 < 16; m590 = m590 + 1) 
        begin: inbit590
            assign data_11[m590 + b590*16 + a21*28*16] = data_11_array[a21][b590][m590];
        end
    endgenerate
    generate 
        localparam integer b591 = 3;
        for (m591 = 0; m591 < 16; m591 = m591 + 1) 
        begin: inbit591
            assign data_11[m591 + b591*16 + a21*28*16] = data_11_array[a21][b591][m591];
        end
    endgenerate
    generate 
        localparam integer b592 = 4;
        for (m592 = 0; m592 < 16; m592 = m592 + 1) 
        begin: inbit592
            assign data_11[m592 + b592*16 + a21*28*16] = data_11_array[a21][b592][m592];
        end
    endgenerate
    generate 
        localparam integer b593 = 5;
        for (m593 = 0; m593 < 16; m593 = m593 + 1) 
        begin: inbit593
            assign data_11[m593 + b593*16 + a21*28*16] = data_11_array[a21][b593][m593];
        end
    endgenerate
    generate 
        localparam integer b594 = 6;
        for (m594 = 0; m594 < 16; m594 = m594 + 1) 
        begin: inbit594
            assign data_11[m594 + b594*16 + a21*28*16] = data_11_array[a21][b594][m594];
        end
    endgenerate
    generate 
        localparam integer b595 = 7;
        for (m595 = 0; m595 < 16; m595 = m595 + 1) 
        begin: inbit595
            assign data_11[m595 + b595*16 + a21*28*16] = data_11_array[a21][b595][m595];
        end
    endgenerate
    generate 
        localparam integer b596 = 8;
        for (m596 = 0; m596 < 16; m596 = m596 + 1) 
        begin: inbit596
            assign data_11[m596 + b596*16 + a21*28*16] = data_11_array[a21][b596][m596];
        end
    endgenerate
    generate 
        localparam integer b597 = 9;
        for (m597 = 0; m597 < 16; m597 = m597 + 1) 
        begin: inbit597
            assign data_11[m597 + b597*16 + a21*28*16] = data_11_array[a21][b597][m597];
        end
    endgenerate
    generate 
        localparam integer b598 = 10;
        for (m598 = 0; m598 < 16; m598 = m598 + 1) 
        begin: inbit598
            assign data_11[m598 + b598*16 + a21*28*16] = data_11_array[a21][b598][m598];
        end
    endgenerate
    generate 
        localparam integer b599 = 11;
        for (m599 = 0; m599 < 16; m599 = m599 + 1) 
        begin: inbit599
            assign data_11[m599 + b599*16 + a21*28*16] = data_11_array[a21][b599][m599];
        end
    endgenerate
    generate 
        localparam integer b600 = 12;
        for (m600 = 0; m600 < 16; m600 = m600 + 1) 
        begin: inbit600
            assign data_11[m600 + b600*16 + a21*28*16] = data_11_array[a21][b600][m600];
        end
    endgenerate
    generate 
        localparam integer b601 = 13;
        for (m601 = 0; m601 < 16; m601 = m601 + 1) 
        begin: inbit601
            assign data_11[m601 + b601*16 + a21*28*16] = data_11_array[a21][b601][m601];
        end
    endgenerate
    generate 
        localparam integer b602 = 14;
        for (m602 = 0; m602 < 16; m602 = m602 + 1) 
        begin: inbit602
            assign data_11[m602 + b602*16 + a21*28*16] = data_11_array[a21][b602][m602];
        end
    endgenerate
    generate 
        localparam integer b603 = 15;
        for (m603 = 0; m603 < 16; m603 = m603 + 1) 
        begin: inbit603
            assign data_11[m603 + b603*16 + a21*28*16] = data_11_array[a21][b603][m603];
        end
    endgenerate
    generate 
        localparam integer b604 = 16;
        for (m604 = 0; m604 < 16; m604 = m604 + 1) 
        begin: inbit604
            assign data_11[m604 + b604*16 + a21*28*16] = data_11_array[a21][b604][m604];
        end
    endgenerate
    generate 
        localparam integer b605 = 17;
        for (m605 = 0; m605 < 16; m605 = m605 + 1) 
        begin: inbit605
            assign data_11[m605 + b605*16 + a21*28*16] = data_11_array[a21][b605][m605];
        end
    endgenerate
    generate 
        localparam integer b606 = 18;
        for (m606 = 0; m606 < 16; m606 = m606 + 1) 
        begin: inbit606
            assign data_11[m606 + b606*16 + a21*28*16] = data_11_array[a21][b606][m606];
        end
    endgenerate
    generate 
        localparam integer b607 = 19;
        for (m607 = 0; m607 < 16; m607 = m607 + 1) 
        begin: inbit607
            assign data_11[m607 + b607*16 + a21*28*16] = data_11_array[a21][b607][m607];
        end
    endgenerate
    generate 
        localparam integer b608 = 20;
        for (m608 = 0; m608 < 16; m608 = m608 + 1) 
        begin: inbit608
            assign data_11[m608 + b608*16 + a21*28*16] = data_11_array[a21][b608][m608];
        end
    endgenerate
    generate 
        localparam integer b609 = 21;
        for (m609 = 0; m609 < 16; m609 = m609 + 1) 
        begin: inbit609
            assign data_11[m609 + b609*16 + a21*28*16] = data_11_array[a21][b609][m609];
        end
    endgenerate
    generate 
        localparam integer b610 = 22;
        for (m610 = 0; m610 < 16; m610 = m610 + 1) 
        begin: inbit610
            assign data_11[m610 + b610*16 + a21*28*16] = data_11_array[a21][b610][m610];
        end
    endgenerate
    generate 
        localparam integer b611 = 23;
        for (m611 = 0; m611 < 16; m611 = m611 + 1) 
        begin: inbit611
            assign data_11[m611 + b611*16 + a21*28*16] = data_11_array[a21][b611][m611];
        end
    endgenerate
    generate 
        localparam integer b612 = 24;
        for (m612 = 0; m612 < 16; m612 = m612 + 1) 
        begin: inbit612
            assign data_11[m612 + b612*16 + a21*28*16] = data_11_array[a21][b612][m612];
        end
    endgenerate
    generate 
        localparam integer b613 = 25;
        for (m613 = 0; m613 < 16; m613 = m613 + 1) 
        begin: inbit613
            assign data_11[m613 + b613*16 + a21*28*16] = data_11_array[a21][b613][m613];
        end
    endgenerate
    generate 
        localparam integer b614 = 26;
        for (m614 = 0; m614 < 16; m614 = m614 + 1) 
        begin: inbit614
            assign data_11[m614 + b614*16 + a21*28*16] = data_11_array[a21][b614][m614];
        end
    endgenerate
    generate 
        localparam integer b615 = 27;
        for (m615 = 0; m615 < 16; m615 = m615 + 1) 
        begin: inbit615
            assign data_11[m615 + b615*16 + a21*28*16] = data_11_array[a21][b615][m615];
        end
    endgenerate
    localparam integer a22 = 22;
    generate 
        localparam integer b616 = 0;
        for (m616 = 0; m616 < 16; m616 = m616 + 1) 
        begin: inbit616
            assign data_11[m616 + b616*16 + a22*28*16] = data_11_array[a22][b616][m616];
        end
    endgenerate
    generate 
        localparam integer b617 = 1;
        for (m617 = 0; m617 < 16; m617 = m617 + 1) 
        begin: inbit617
            assign data_11[m617 + b617*16 + a22*28*16] = data_11_array[a22][b617][m617];
        end
    endgenerate
    generate 
        localparam integer b618 = 2;
        for (m618 = 0; m618 < 16; m618 = m618 + 1) 
        begin: inbit618
            assign data_11[m618 + b618*16 + a22*28*16] = data_11_array[a22][b618][m618];
        end
    endgenerate
    generate 
        localparam integer b619 = 3;
        for (m619 = 0; m619 < 16; m619 = m619 + 1) 
        begin: inbit619
            assign data_11[m619 + b619*16 + a22*28*16] = data_11_array[a22][b619][m619];
        end
    endgenerate
    generate 
        localparam integer b620 = 4;
        for (m620 = 0; m620 < 16; m620 = m620 + 1) 
        begin: inbit620
            assign data_11[m620 + b620*16 + a22*28*16] = data_11_array[a22][b620][m620];
        end
    endgenerate
    generate 
        localparam integer b621 = 5;
        for (m621 = 0; m621 < 16; m621 = m621 + 1) 
        begin: inbit621
            assign data_11[m621 + b621*16 + a22*28*16] = data_11_array[a22][b621][m621];
        end
    endgenerate
    generate 
        localparam integer b622 = 6;
        for (m622 = 0; m622 < 16; m622 = m622 + 1) 
        begin: inbit622
            assign data_11[m622 + b622*16 + a22*28*16] = data_11_array[a22][b622][m622];
        end
    endgenerate
    generate 
        localparam integer b623 = 7;
        for (m623 = 0; m623 < 16; m623 = m623 + 1) 
        begin: inbit623
            assign data_11[m623 + b623*16 + a22*28*16] = data_11_array[a22][b623][m623];
        end
    endgenerate
    generate 
        localparam integer b624 = 8;
        for (m624 = 0; m624 < 16; m624 = m624 + 1) 
        begin: inbit624
            assign data_11[m624 + b624*16 + a22*28*16] = data_11_array[a22][b624][m624];
        end
    endgenerate
    generate 
        localparam integer b625 = 9;
        for (m625 = 0; m625 < 16; m625 = m625 + 1) 
        begin: inbit625
            assign data_11[m625 + b625*16 + a22*28*16] = data_11_array[a22][b625][m625];
        end
    endgenerate
    generate 
        localparam integer b626 = 10;
        for (m626 = 0; m626 < 16; m626 = m626 + 1) 
        begin: inbit626
            assign data_11[m626 + b626*16 + a22*28*16] = data_11_array[a22][b626][m626];
        end
    endgenerate
    generate 
        localparam integer b627 = 11;
        for (m627 = 0; m627 < 16; m627 = m627 + 1) 
        begin: inbit627
            assign data_11[m627 + b627*16 + a22*28*16] = data_11_array[a22][b627][m627];
        end
    endgenerate
    generate 
        localparam integer b628 = 12;
        for (m628 = 0; m628 < 16; m628 = m628 + 1) 
        begin: inbit628
            assign data_11[m628 + b628*16 + a22*28*16] = data_11_array[a22][b628][m628];
        end
    endgenerate
    generate 
        localparam integer b629 = 13;
        for (m629 = 0; m629 < 16; m629 = m629 + 1) 
        begin: inbit629
            assign data_11[m629 + b629*16 + a22*28*16] = data_11_array[a22][b629][m629];
        end
    endgenerate
    generate 
        localparam integer b630 = 14;
        for (m630 = 0; m630 < 16; m630 = m630 + 1) 
        begin: inbit630
            assign data_11[m630 + b630*16 + a22*28*16] = data_11_array[a22][b630][m630];
        end
    endgenerate
    generate 
        localparam integer b631 = 15;
        for (m631 = 0; m631 < 16; m631 = m631 + 1) 
        begin: inbit631
            assign data_11[m631 + b631*16 + a22*28*16] = data_11_array[a22][b631][m631];
        end
    endgenerate
    generate 
        localparam integer b632 = 16;
        for (m632 = 0; m632 < 16; m632 = m632 + 1) 
        begin: inbit632
            assign data_11[m632 + b632*16 + a22*28*16] = data_11_array[a22][b632][m632];
        end
    endgenerate
    generate 
        localparam integer b633 = 17;
        for (m633 = 0; m633 < 16; m633 = m633 + 1) 
        begin: inbit633
            assign data_11[m633 + b633*16 + a22*28*16] = data_11_array[a22][b633][m633];
        end
    endgenerate
    generate 
        localparam integer b634 = 18;
        for (m634 = 0; m634 < 16; m634 = m634 + 1) 
        begin: inbit634
            assign data_11[m634 + b634*16 + a22*28*16] = data_11_array[a22][b634][m634];
        end
    endgenerate
    generate 
        localparam integer b635 = 19;
        for (m635 = 0; m635 < 16; m635 = m635 + 1) 
        begin: inbit635
            assign data_11[m635 + b635*16 + a22*28*16] = data_11_array[a22][b635][m635];
        end
    endgenerate
    generate 
        localparam integer b636 = 20;
        for (m636 = 0; m636 < 16; m636 = m636 + 1) 
        begin: inbit636
            assign data_11[m636 + b636*16 + a22*28*16] = data_11_array[a22][b636][m636];
        end
    endgenerate
    generate 
        localparam integer b637 = 21;
        for (m637 = 0; m637 < 16; m637 = m637 + 1) 
        begin: inbit637
            assign data_11[m637 + b637*16 + a22*28*16] = data_11_array[a22][b637][m637];
        end
    endgenerate
    generate 
        localparam integer b638 = 22;
        for (m638 = 0; m638 < 16; m638 = m638 + 1) 
        begin: inbit638
            assign data_11[m638 + b638*16 + a22*28*16] = data_11_array[a22][b638][m638];
        end
    endgenerate
    generate 
        localparam integer b639 = 23;
        for (m639 = 0; m639 < 16; m639 = m639 + 1) 
        begin: inbit639
            assign data_11[m639 + b639*16 + a22*28*16] = data_11_array[a22][b639][m639];
        end
    endgenerate
    generate 
        localparam integer b640 = 24;
        for (m640 = 0; m640 < 16; m640 = m640 + 1) 
        begin: inbit640
            assign data_11[m640 + b640*16 + a22*28*16] = data_11_array[a22][b640][m640];
        end
    endgenerate
    generate 
        localparam integer b641 = 25;
        for (m641 = 0; m641 < 16; m641 = m641 + 1) 
        begin: inbit641
            assign data_11[m641 + b641*16 + a22*28*16] = data_11_array[a22][b641][m641];
        end
    endgenerate
    generate 
        localparam integer b642 = 26;
        for (m642 = 0; m642 < 16; m642 = m642 + 1) 
        begin: inbit642
            assign data_11[m642 + b642*16 + a22*28*16] = data_11_array[a22][b642][m642];
        end
    endgenerate
    generate 
        localparam integer b643 = 27;
        for (m643 = 0; m643 < 16; m643 = m643 + 1) 
        begin: inbit643
            assign data_11[m643 + b643*16 + a22*28*16] = data_11_array[a22][b643][m643];
        end
    endgenerate
    localparam integer a23 = 23;
    generate 
        localparam integer b644 = 0;
        for (m644 = 0; m644 < 16; m644 = m644 + 1) 
        begin: inbit644
            assign data_11[m644 + b644*16 + a23*28*16] = data_11_array[a23][b644][m644];
        end
    endgenerate
    generate 
        localparam integer b645 = 1;
        for (m645 = 0; m645 < 16; m645 = m645 + 1) 
        begin: inbit645
            assign data_11[m645 + b645*16 + a23*28*16] = data_11_array[a23][b645][m645];
        end
    endgenerate
    generate 
        localparam integer b646 = 2;
        for (m646 = 0; m646 < 16; m646 = m646 + 1) 
        begin: inbit646
            assign data_11[m646 + b646*16 + a23*28*16] = data_11_array[a23][b646][m646];
        end
    endgenerate
    generate 
        localparam integer b647 = 3;
        for (m647 = 0; m647 < 16; m647 = m647 + 1) 
        begin: inbit647
            assign data_11[m647 + b647*16 + a23*28*16] = data_11_array[a23][b647][m647];
        end
    endgenerate
    generate 
        localparam integer b648 = 4;
        for (m648 = 0; m648 < 16; m648 = m648 + 1) 
        begin: inbit648
            assign data_11[m648 + b648*16 + a23*28*16] = data_11_array[a23][b648][m648];
        end
    endgenerate
    generate 
        localparam integer b649 = 5;
        for (m649 = 0; m649 < 16; m649 = m649 + 1) 
        begin: inbit649
            assign data_11[m649 + b649*16 + a23*28*16] = data_11_array[a23][b649][m649];
        end
    endgenerate
    generate 
        localparam integer b650 = 6;
        for (m650 = 0; m650 < 16; m650 = m650 + 1) 
        begin: inbit650
            assign data_11[m650 + b650*16 + a23*28*16] = data_11_array[a23][b650][m650];
        end
    endgenerate
    generate 
        localparam integer b651 = 7;
        for (m651 = 0; m651 < 16; m651 = m651 + 1) 
        begin: inbit651
            assign data_11[m651 + b651*16 + a23*28*16] = data_11_array[a23][b651][m651];
        end
    endgenerate
    generate 
        localparam integer b652 = 8;
        for (m652 = 0; m652 < 16; m652 = m652 + 1) 
        begin: inbit652
            assign data_11[m652 + b652*16 + a23*28*16] = data_11_array[a23][b652][m652];
        end
    endgenerate
    generate 
        localparam integer b653 = 9;
        for (m653 = 0; m653 < 16; m653 = m653 + 1) 
        begin: inbit653
            assign data_11[m653 + b653*16 + a23*28*16] = data_11_array[a23][b653][m653];
        end
    endgenerate
    generate 
        localparam integer b654 = 10;
        for (m654 = 0; m654 < 16; m654 = m654 + 1) 
        begin: inbit654
            assign data_11[m654 + b654*16 + a23*28*16] = data_11_array[a23][b654][m654];
        end
    endgenerate
    generate 
        localparam integer b655 = 11;
        for (m655 = 0; m655 < 16; m655 = m655 + 1) 
        begin: inbit655
            assign data_11[m655 + b655*16 + a23*28*16] = data_11_array[a23][b655][m655];
        end
    endgenerate
    generate 
        localparam integer b656 = 12;
        for (m656 = 0; m656 < 16; m656 = m656 + 1) 
        begin: inbit656
            assign data_11[m656 + b656*16 + a23*28*16] = data_11_array[a23][b656][m656];
        end
    endgenerate
    generate 
        localparam integer b657 = 13;
        for (m657 = 0; m657 < 16; m657 = m657 + 1) 
        begin: inbit657
            assign data_11[m657 + b657*16 + a23*28*16] = data_11_array[a23][b657][m657];
        end
    endgenerate
    generate 
        localparam integer b658 = 14;
        for (m658 = 0; m658 < 16; m658 = m658 + 1) 
        begin: inbit658
            assign data_11[m658 + b658*16 + a23*28*16] = data_11_array[a23][b658][m658];
        end
    endgenerate
    generate 
        localparam integer b659 = 15;
        for (m659 = 0; m659 < 16; m659 = m659 + 1) 
        begin: inbit659
            assign data_11[m659 + b659*16 + a23*28*16] = data_11_array[a23][b659][m659];
        end
    endgenerate
    generate 
        localparam integer b660 = 16;
        for (m660 = 0; m660 < 16; m660 = m660 + 1) 
        begin: inbit660
            assign data_11[m660 + b660*16 + a23*28*16] = data_11_array[a23][b660][m660];
        end
    endgenerate
    generate 
        localparam integer b661 = 17;
        for (m661 = 0; m661 < 16; m661 = m661 + 1) 
        begin: inbit661
            assign data_11[m661 + b661*16 + a23*28*16] = data_11_array[a23][b661][m661];
        end
    endgenerate
    generate 
        localparam integer b662 = 18;
        for (m662 = 0; m662 < 16; m662 = m662 + 1) 
        begin: inbit662
            assign data_11[m662 + b662*16 + a23*28*16] = data_11_array[a23][b662][m662];
        end
    endgenerate
    generate 
        localparam integer b663 = 19;
        for (m663 = 0; m663 < 16; m663 = m663 + 1) 
        begin: inbit663
            assign data_11[m663 + b663*16 + a23*28*16] = data_11_array[a23][b663][m663];
        end
    endgenerate
    generate 
        localparam integer b664 = 20;
        for (m664 = 0; m664 < 16; m664 = m664 + 1) 
        begin: inbit664
            assign data_11[m664 + b664*16 + a23*28*16] = data_11_array[a23][b664][m664];
        end
    endgenerate
    generate 
        localparam integer b665 = 21;
        for (m665 = 0; m665 < 16; m665 = m665 + 1) 
        begin: inbit665
            assign data_11[m665 + b665*16 + a23*28*16] = data_11_array[a23][b665][m665];
        end
    endgenerate
    generate 
        localparam integer b666 = 22;
        for (m666 = 0; m666 < 16; m666 = m666 + 1) 
        begin: inbit666
            assign data_11[m666 + b666*16 + a23*28*16] = data_11_array[a23][b666][m666];
        end
    endgenerate
    generate 
        localparam integer b667 = 23;
        for (m667 = 0; m667 < 16; m667 = m667 + 1) 
        begin: inbit667
            assign data_11[m667 + b667*16 + a23*28*16] = data_11_array[a23][b667][m667];
        end
    endgenerate
    generate 
        localparam integer b668 = 24;
        for (m668 = 0; m668 < 16; m668 = m668 + 1) 
        begin: inbit668
            assign data_11[m668 + b668*16 + a23*28*16] = data_11_array[a23][b668][m668];
        end
    endgenerate
    generate 
        localparam integer b669 = 25;
        for (m669 = 0; m669 < 16; m669 = m669 + 1) 
        begin: inbit669
            assign data_11[m669 + b669*16 + a23*28*16] = data_11_array[a23][b669][m669];
        end
    endgenerate
    generate 
        localparam integer b670 = 26;
        for (m670 = 0; m670 < 16; m670 = m670 + 1) 
        begin: inbit670
            assign data_11[m670 + b670*16 + a23*28*16] = data_11_array[a23][b670][m670];
        end
    endgenerate
    generate 
        localparam integer b671 = 27;
        for (m671 = 0; m671 < 16; m671 = m671 + 1) 
        begin: inbit671
            assign data_11[m671 + b671*16 + a23*28*16] = data_11_array[a23][b671][m671];
        end
    endgenerate
    localparam integer a24 = 24;
    generate 
        localparam integer b672 = 0;
        for (m672 = 0; m672 < 16; m672 = m672 + 1) 
        begin: inbit672
            assign data_11[m672 + b672*16 + a24*28*16] = data_11_array[a24][b672][m672];
        end
    endgenerate
    generate 
        localparam integer b673 = 1;
        for (m673 = 0; m673 < 16; m673 = m673 + 1) 
        begin: inbit673
            assign data_11[m673 + b673*16 + a24*28*16] = data_11_array[a24][b673][m673];
        end
    endgenerate
    generate 
        localparam integer b674 = 2;
        for (m674 = 0; m674 < 16; m674 = m674 + 1) 
        begin: inbit674
            assign data_11[m674 + b674*16 + a24*28*16] = data_11_array[a24][b674][m674];
        end
    endgenerate
    generate 
        localparam integer b675 = 3;
        for (m675 = 0; m675 < 16; m675 = m675 + 1) 
        begin: inbit675
            assign data_11[m675 + b675*16 + a24*28*16] = data_11_array[a24][b675][m675];
        end
    endgenerate
    generate 
        localparam integer b676 = 4;
        for (m676 = 0; m676 < 16; m676 = m676 + 1) 
        begin: inbit676
            assign data_11[m676 + b676*16 + a24*28*16] = data_11_array[a24][b676][m676];
        end
    endgenerate
    generate 
        localparam integer b677 = 5;
        for (m677 = 0; m677 < 16; m677 = m677 + 1) 
        begin: inbit677
            assign data_11[m677 + b677*16 + a24*28*16] = data_11_array[a24][b677][m677];
        end
    endgenerate
    generate 
        localparam integer b678 = 6;
        for (m678 = 0; m678 < 16; m678 = m678 + 1) 
        begin: inbit678
            assign data_11[m678 + b678*16 + a24*28*16] = data_11_array[a24][b678][m678];
        end
    endgenerate
    generate 
        localparam integer b679 = 7;
        for (m679 = 0; m679 < 16; m679 = m679 + 1) 
        begin: inbit679
            assign data_11[m679 + b679*16 + a24*28*16] = data_11_array[a24][b679][m679];
        end
    endgenerate
    generate 
        localparam integer b680 = 8;
        for (m680 = 0; m680 < 16; m680 = m680 + 1) 
        begin: inbit680
            assign data_11[m680 + b680*16 + a24*28*16] = data_11_array[a24][b680][m680];
        end
    endgenerate
    generate 
        localparam integer b681 = 9;
        for (m681 = 0; m681 < 16; m681 = m681 + 1) 
        begin: inbit681
            assign data_11[m681 + b681*16 + a24*28*16] = data_11_array[a24][b681][m681];
        end
    endgenerate
    generate 
        localparam integer b682 = 10;
        for (m682 = 0; m682 < 16; m682 = m682 + 1) 
        begin: inbit682
            assign data_11[m682 + b682*16 + a24*28*16] = data_11_array[a24][b682][m682];
        end
    endgenerate
    generate 
        localparam integer b683 = 11;
        for (m683 = 0; m683 < 16; m683 = m683 + 1) 
        begin: inbit683
            assign data_11[m683 + b683*16 + a24*28*16] = data_11_array[a24][b683][m683];
        end
    endgenerate
    generate 
        localparam integer b684 = 12;
        for (m684 = 0; m684 < 16; m684 = m684 + 1) 
        begin: inbit684
            assign data_11[m684 + b684*16 + a24*28*16] = data_11_array[a24][b684][m684];
        end
    endgenerate
    generate 
        localparam integer b685 = 13;
        for (m685 = 0; m685 < 16; m685 = m685 + 1) 
        begin: inbit685
            assign data_11[m685 + b685*16 + a24*28*16] = data_11_array[a24][b685][m685];
        end
    endgenerate
    generate 
        localparam integer b686 = 14;
        for (m686 = 0; m686 < 16; m686 = m686 + 1) 
        begin: inbit686
            assign data_11[m686 + b686*16 + a24*28*16] = data_11_array[a24][b686][m686];
        end
    endgenerate
    generate 
        localparam integer b687 = 15;
        for (m687 = 0; m687 < 16; m687 = m687 + 1) 
        begin: inbit687
            assign data_11[m687 + b687*16 + a24*28*16] = data_11_array[a24][b687][m687];
        end
    endgenerate
    generate 
        localparam integer b688 = 16;
        for (m688 = 0; m688 < 16; m688 = m688 + 1) 
        begin: inbit688
            assign data_11[m688 + b688*16 + a24*28*16] = data_11_array[a24][b688][m688];
        end
    endgenerate
    generate 
        localparam integer b689 = 17;
        for (m689 = 0; m689 < 16; m689 = m689 + 1) 
        begin: inbit689
            assign data_11[m689 + b689*16 + a24*28*16] = data_11_array[a24][b689][m689];
        end
    endgenerate
    generate 
        localparam integer b690 = 18;
        for (m690 = 0; m690 < 16; m690 = m690 + 1) 
        begin: inbit690
            assign data_11[m690 + b690*16 + a24*28*16] = data_11_array[a24][b690][m690];
        end
    endgenerate
    generate 
        localparam integer b691 = 19;
        for (m691 = 0; m691 < 16; m691 = m691 + 1) 
        begin: inbit691
            assign data_11[m691 + b691*16 + a24*28*16] = data_11_array[a24][b691][m691];
        end
    endgenerate
    generate 
        localparam integer b692 = 20;
        for (m692 = 0; m692 < 16; m692 = m692 + 1) 
        begin: inbit692
            assign data_11[m692 + b692*16 + a24*28*16] = data_11_array[a24][b692][m692];
        end
    endgenerate
    generate 
        localparam integer b693 = 21;
        for (m693 = 0; m693 < 16; m693 = m693 + 1) 
        begin: inbit693
            assign data_11[m693 + b693*16 + a24*28*16] = data_11_array[a24][b693][m693];
        end
    endgenerate
    generate 
        localparam integer b694 = 22;
        for (m694 = 0; m694 < 16; m694 = m694 + 1) 
        begin: inbit694
            assign data_11[m694 + b694*16 + a24*28*16] = data_11_array[a24][b694][m694];
        end
    endgenerate
    generate 
        localparam integer b695 = 23;
        for (m695 = 0; m695 < 16; m695 = m695 + 1) 
        begin: inbit695
            assign data_11[m695 + b695*16 + a24*28*16] = data_11_array[a24][b695][m695];
        end
    endgenerate
    generate 
        localparam integer b696 = 24;
        for (m696 = 0; m696 < 16; m696 = m696 + 1) 
        begin: inbit696
            assign data_11[m696 + b696*16 + a24*28*16] = data_11_array[a24][b696][m696];
        end
    endgenerate
    generate 
        localparam integer b697 = 25;
        for (m697 = 0; m697 < 16; m697 = m697 + 1) 
        begin: inbit697
            assign data_11[m697 + b697*16 + a24*28*16] = data_11_array[a24][b697][m697];
        end
    endgenerate
    generate 
        localparam integer b698 = 26;
        for (m698 = 0; m698 < 16; m698 = m698 + 1) 
        begin: inbit698
            assign data_11[m698 + b698*16 + a24*28*16] = data_11_array[a24][b698][m698];
        end
    endgenerate
    generate 
        localparam integer b699 = 27;
        for (m699 = 0; m699 < 16; m699 = m699 + 1) 
        begin: inbit699
            assign data_11[m699 + b699*16 + a24*28*16] = data_11_array[a24][b699][m699];
        end
    endgenerate
    localparam integer a25 = 25;
    generate 
        localparam integer b700 = 0;
        for (m700 = 0; m700 < 16; m700 = m700 + 1) 
        begin: inbit700
            assign data_11[m700 + b700*16 + a25*28*16] = data_11_array[a25][b700][m700];
        end
    endgenerate
    generate 
        localparam integer b701 = 1;
        for (m701 = 0; m701 < 16; m701 = m701 + 1) 
        begin: inbit701
            assign data_11[m701 + b701*16 + a25*28*16] = data_11_array[a25][b701][m701];
        end
    endgenerate
    generate 
        localparam integer b702 = 2;
        for (m702 = 0; m702 < 16; m702 = m702 + 1) 
        begin: inbit702
            assign data_11[m702 + b702*16 + a25*28*16] = data_11_array[a25][b702][m702];
        end
    endgenerate
    generate 
        localparam integer b703 = 3;
        for (m703 = 0; m703 < 16; m703 = m703 + 1) 
        begin: inbit703
            assign data_11[m703 + b703*16 + a25*28*16] = data_11_array[a25][b703][m703];
        end
    endgenerate
    generate 
        localparam integer b704 = 4;
        for (m704 = 0; m704 < 16; m704 = m704 + 1) 
        begin: inbit704
            assign data_11[m704 + b704*16 + a25*28*16] = data_11_array[a25][b704][m704];
        end
    endgenerate
    generate 
        localparam integer b705 = 5;
        for (m705 = 0; m705 < 16; m705 = m705 + 1) 
        begin: inbit705
            assign data_11[m705 + b705*16 + a25*28*16] = data_11_array[a25][b705][m705];
        end
    endgenerate
    generate 
        localparam integer b706 = 6;
        for (m706 = 0; m706 < 16; m706 = m706 + 1) 
        begin: inbit706
            assign data_11[m706 + b706*16 + a25*28*16] = data_11_array[a25][b706][m706];
        end
    endgenerate
    generate 
        localparam integer b707 = 7;
        for (m707 = 0; m707 < 16; m707 = m707 + 1) 
        begin: inbit707
            assign data_11[m707 + b707*16 + a25*28*16] = data_11_array[a25][b707][m707];
        end
    endgenerate
    generate 
        localparam integer b708 = 8;
        for (m708 = 0; m708 < 16; m708 = m708 + 1) 
        begin: inbit708
            assign data_11[m708 + b708*16 + a25*28*16] = data_11_array[a25][b708][m708];
        end
    endgenerate
    generate 
        localparam integer b709 = 9;
        for (m709 = 0; m709 < 16; m709 = m709 + 1) 
        begin: inbit709
            assign data_11[m709 + b709*16 + a25*28*16] = data_11_array[a25][b709][m709];
        end
    endgenerate
    generate 
        localparam integer b710 = 10;
        for (m710 = 0; m710 < 16; m710 = m710 + 1) 
        begin: inbit710
            assign data_11[m710 + b710*16 + a25*28*16] = data_11_array[a25][b710][m710];
        end
    endgenerate
    generate 
        localparam integer b711 = 11;
        for (m711 = 0; m711 < 16; m711 = m711 + 1) 
        begin: inbit711
            assign data_11[m711 + b711*16 + a25*28*16] = data_11_array[a25][b711][m711];
        end
    endgenerate
    generate 
        localparam integer b712 = 12;
        for (m712 = 0; m712 < 16; m712 = m712 + 1) 
        begin: inbit712
            assign data_11[m712 + b712*16 + a25*28*16] = data_11_array[a25][b712][m712];
        end
    endgenerate
    generate 
        localparam integer b713 = 13;
        for (m713 = 0; m713 < 16; m713 = m713 + 1) 
        begin: inbit713
            assign data_11[m713 + b713*16 + a25*28*16] = data_11_array[a25][b713][m713];
        end
    endgenerate
    generate 
        localparam integer b714 = 14;
        for (m714 = 0; m714 < 16; m714 = m714 + 1) 
        begin: inbit714
            assign data_11[m714 + b714*16 + a25*28*16] = data_11_array[a25][b714][m714];
        end
    endgenerate
    generate 
        localparam integer b715 = 15;
        for (m715 = 0; m715 < 16; m715 = m715 + 1) 
        begin: inbit715
            assign data_11[m715 + b715*16 + a25*28*16] = data_11_array[a25][b715][m715];
        end
    endgenerate
    generate 
        localparam integer b716 = 16;
        for (m716 = 0; m716 < 16; m716 = m716 + 1) 
        begin: inbit716
            assign data_11[m716 + b716*16 + a25*28*16] = data_11_array[a25][b716][m716];
        end
    endgenerate
    generate 
        localparam integer b717 = 17;
        for (m717 = 0; m717 < 16; m717 = m717 + 1) 
        begin: inbit717
            assign data_11[m717 + b717*16 + a25*28*16] = data_11_array[a25][b717][m717];
        end
    endgenerate
    generate 
        localparam integer b718 = 18;
        for (m718 = 0; m718 < 16; m718 = m718 + 1) 
        begin: inbit718
            assign data_11[m718 + b718*16 + a25*28*16] = data_11_array[a25][b718][m718];
        end
    endgenerate
    generate 
        localparam integer b719 = 19;
        for (m719 = 0; m719 < 16; m719 = m719 + 1) 
        begin: inbit719
            assign data_11[m719 + b719*16 + a25*28*16] = data_11_array[a25][b719][m719];
        end
    endgenerate
    generate 
        localparam integer b720 = 20;
        for (m720 = 0; m720 < 16; m720 = m720 + 1) 
        begin: inbit720
            assign data_11[m720 + b720*16 + a25*28*16] = data_11_array[a25][b720][m720];
        end
    endgenerate
    generate 
        localparam integer b721 = 21;
        for (m721 = 0; m721 < 16; m721 = m721 + 1) 
        begin: inbit721
            assign data_11[m721 + b721*16 + a25*28*16] = data_11_array[a25][b721][m721];
        end
    endgenerate
    generate 
        localparam integer b722 = 22;
        for (m722 = 0; m722 < 16; m722 = m722 + 1) 
        begin: inbit722
            assign data_11[m722 + b722*16 + a25*28*16] = data_11_array[a25][b722][m722];
        end
    endgenerate
    generate 
        localparam integer b723 = 23;
        for (m723 = 0; m723 < 16; m723 = m723 + 1) 
        begin: inbit723
            assign data_11[m723 + b723*16 + a25*28*16] = data_11_array[a25][b723][m723];
        end
    endgenerate
    generate 
        localparam integer b724 = 24;
        for (m724 = 0; m724 < 16; m724 = m724 + 1) 
        begin: inbit724
            assign data_11[m724 + b724*16 + a25*28*16] = data_11_array[a25][b724][m724];
        end
    endgenerate
    generate 
        localparam integer b725 = 25;
        for (m725 = 0; m725 < 16; m725 = m725 + 1) 
        begin: inbit725
            assign data_11[m725 + b725*16 + a25*28*16] = data_11_array[a25][b725][m725];
        end
    endgenerate
    generate 
        localparam integer b726 = 26;
        for (m726 = 0; m726 < 16; m726 = m726 + 1) 
        begin: inbit726
            assign data_11[m726 + b726*16 + a25*28*16] = data_11_array[a25][b726][m726];
        end
    endgenerate
    generate 
        localparam integer b727 = 27;
        for (m727 = 0; m727 < 16; m727 = m727 + 1) 
        begin: inbit727
            assign data_11[m727 + b727*16 + a25*28*16] = data_11_array[a25][b727][m727];
        end
    endgenerate
    localparam integer a26 = 26;
    generate 
        localparam integer b728 = 0;
        for (m728 = 0; m728 < 16; m728 = m728 + 1) 
        begin: inbit728
            assign data_11[m728 + b728*16 + a26*28*16] = data_11_array[a26][b728][m728];
        end
    endgenerate
    generate 
        localparam integer b729 = 1;
        for (m729 = 0; m729 < 16; m729 = m729 + 1) 
        begin: inbit729
            assign data_11[m729 + b729*16 + a26*28*16] = data_11_array[a26][b729][m729];
        end
    endgenerate
    generate 
        localparam integer b730 = 2;
        for (m730 = 0; m730 < 16; m730 = m730 + 1) 
        begin: inbit730
            assign data_11[m730 + b730*16 + a26*28*16] = data_11_array[a26][b730][m730];
        end
    endgenerate
    generate 
        localparam integer b731 = 3;
        for (m731 = 0; m731 < 16; m731 = m731 + 1) 
        begin: inbit731
            assign data_11[m731 + b731*16 + a26*28*16] = data_11_array[a26][b731][m731];
        end
    endgenerate
    generate 
        localparam integer b732 = 4;
        for (m732 = 0; m732 < 16; m732 = m732 + 1) 
        begin: inbit732
            assign data_11[m732 + b732*16 + a26*28*16] = data_11_array[a26][b732][m732];
        end
    endgenerate
    generate 
        localparam integer b733 = 5;
        for (m733 = 0; m733 < 16; m733 = m733 + 1) 
        begin: inbit733
            assign data_11[m733 + b733*16 + a26*28*16] = data_11_array[a26][b733][m733];
        end
    endgenerate
    generate 
        localparam integer b734 = 6;
        for (m734 = 0; m734 < 16; m734 = m734 + 1) 
        begin: inbit734
            assign data_11[m734 + b734*16 + a26*28*16] = data_11_array[a26][b734][m734];
        end
    endgenerate
    generate 
        localparam integer b735 = 7;
        for (m735 = 0; m735 < 16; m735 = m735 + 1) 
        begin: inbit735
            assign data_11[m735 + b735*16 + a26*28*16] = data_11_array[a26][b735][m735];
        end
    endgenerate
    generate 
        localparam integer b736 = 8;
        for (m736 = 0; m736 < 16; m736 = m736 + 1) 
        begin: inbit736
            assign data_11[m736 + b736*16 + a26*28*16] = data_11_array[a26][b736][m736];
        end
    endgenerate
    generate 
        localparam integer b737 = 9;
        for (m737 = 0; m737 < 16; m737 = m737 + 1) 
        begin: inbit737
            assign data_11[m737 + b737*16 + a26*28*16] = data_11_array[a26][b737][m737];
        end
    endgenerate
    generate 
        localparam integer b738 = 10;
        for (m738 = 0; m738 < 16; m738 = m738 + 1) 
        begin: inbit738
            assign data_11[m738 + b738*16 + a26*28*16] = data_11_array[a26][b738][m738];
        end
    endgenerate
    generate 
        localparam integer b739 = 11;
        for (m739 = 0; m739 < 16; m739 = m739 + 1) 
        begin: inbit739
            assign data_11[m739 + b739*16 + a26*28*16] = data_11_array[a26][b739][m739];
        end
    endgenerate
    generate 
        localparam integer b740 = 12;
        for (m740 = 0; m740 < 16; m740 = m740 + 1) 
        begin: inbit740
            assign data_11[m740 + b740*16 + a26*28*16] = data_11_array[a26][b740][m740];
        end
    endgenerate
    generate 
        localparam integer b741 = 13;
        for (m741 = 0; m741 < 16; m741 = m741 + 1) 
        begin: inbit741
            assign data_11[m741 + b741*16 + a26*28*16] = data_11_array[a26][b741][m741];
        end
    endgenerate
    generate 
        localparam integer b742 = 14;
        for (m742 = 0; m742 < 16; m742 = m742 + 1) 
        begin: inbit742
            assign data_11[m742 + b742*16 + a26*28*16] = data_11_array[a26][b742][m742];
        end
    endgenerate
    generate 
        localparam integer b743 = 15;
        for (m743 = 0; m743 < 16; m743 = m743 + 1) 
        begin: inbit743
            assign data_11[m743 + b743*16 + a26*28*16] = data_11_array[a26][b743][m743];
        end
    endgenerate
    generate 
        localparam integer b744 = 16;
        for (m744 = 0; m744 < 16; m744 = m744 + 1) 
        begin: inbit744
            assign data_11[m744 + b744*16 + a26*28*16] = data_11_array[a26][b744][m744];
        end
    endgenerate
    generate 
        localparam integer b745 = 17;
        for (m745 = 0; m745 < 16; m745 = m745 + 1) 
        begin: inbit745
            assign data_11[m745 + b745*16 + a26*28*16] = data_11_array[a26][b745][m745];
        end
    endgenerate
    generate 
        localparam integer b746 = 18;
        for (m746 = 0; m746 < 16; m746 = m746 + 1) 
        begin: inbit746
            assign data_11[m746 + b746*16 + a26*28*16] = data_11_array[a26][b746][m746];
        end
    endgenerate
    generate 
        localparam integer b747 = 19;
        for (m747 = 0; m747 < 16; m747 = m747 + 1) 
        begin: inbit747
            assign data_11[m747 + b747*16 + a26*28*16] = data_11_array[a26][b747][m747];
        end
    endgenerate
    generate 
        localparam integer b748 = 20;
        for (m748 = 0; m748 < 16; m748 = m748 + 1) 
        begin: inbit748
            assign data_11[m748 + b748*16 + a26*28*16] = data_11_array[a26][b748][m748];
        end
    endgenerate
    generate 
        localparam integer b749 = 21;
        for (m749 = 0; m749 < 16; m749 = m749 + 1) 
        begin: inbit749
            assign data_11[m749 + b749*16 + a26*28*16] = data_11_array[a26][b749][m749];
        end
    endgenerate
    generate 
        localparam integer b750 = 22;
        for (m750 = 0; m750 < 16; m750 = m750 + 1) 
        begin: inbit750
            assign data_11[m750 + b750*16 + a26*28*16] = data_11_array[a26][b750][m750];
        end
    endgenerate
    generate 
        localparam integer b751 = 23;
        for (m751 = 0; m751 < 16; m751 = m751 + 1) 
        begin: inbit751
            assign data_11[m751 + b751*16 + a26*28*16] = data_11_array[a26][b751][m751];
        end
    endgenerate
    generate 
        localparam integer b752 = 24;
        for (m752 = 0; m752 < 16; m752 = m752 + 1) 
        begin: inbit752
            assign data_11[m752 + b752*16 + a26*28*16] = data_11_array[a26][b752][m752];
        end
    endgenerate
    generate 
        localparam integer b753 = 25;
        for (m753 = 0; m753 < 16; m753 = m753 + 1) 
        begin: inbit753
            assign data_11[m753 + b753*16 + a26*28*16] = data_11_array[a26][b753][m753];
        end
    endgenerate
    generate 
        localparam integer b754 = 26;
        for (m754 = 0; m754 < 16; m754 = m754 + 1) 
        begin: inbit754
            assign data_11[m754 + b754*16 + a26*28*16] = data_11_array[a26][b754][m754];
        end
    endgenerate
    generate 
        localparam integer b755 = 27;
        for (m755 = 0; m755 < 16; m755 = m755 + 1) 
        begin: inbit755
            assign data_11[m755 + b755*16 + a26*28*16] = data_11_array[a26][b755][m755];
        end
    endgenerate
    localparam integer a27 = 27;
    generate 
        localparam integer b756 = 0;
        for (m756 = 0; m756 < 16; m756 = m756 + 1) 
        begin: inbit756
            assign data_11[m756 + b756*16 + a27*28*16] = data_11_array[a27][b756][m756];
        end
    endgenerate
    generate 
        localparam integer b757 = 1;
        for (m757 = 0; m757 < 16; m757 = m757 + 1) 
        begin: inbit757
            assign data_11[m757 + b757*16 + a27*28*16] = data_11_array[a27][b757][m757];
        end
    endgenerate
    generate 
        localparam integer b758 = 2;
        for (m758 = 0; m758 < 16; m758 = m758 + 1) 
        begin: inbit758
            assign data_11[m758 + b758*16 + a27*28*16] = data_11_array[a27][b758][m758];
        end
    endgenerate
    generate 
        localparam integer b759 = 3;
        for (m759 = 0; m759 < 16; m759 = m759 + 1) 
        begin: inbit759
            assign data_11[m759 + b759*16 + a27*28*16] = data_11_array[a27][b759][m759];
        end
    endgenerate
    generate 
        localparam integer b760 = 4;
        for (m760 = 0; m760 < 16; m760 = m760 + 1) 
        begin: inbit760
            assign data_11[m760 + b760*16 + a27*28*16] = data_11_array[a27][b760][m760];
        end
    endgenerate
    generate 
        localparam integer b761 = 5;
        for (m761 = 0; m761 < 16; m761 = m761 + 1) 
        begin: inbit761
            assign data_11[m761 + b761*16 + a27*28*16] = data_11_array[a27][b761][m761];
        end
    endgenerate
    generate 
        localparam integer b762 = 6;
        for (m762 = 0; m762 < 16; m762 = m762 + 1) 
        begin: inbit762
            assign data_11[m762 + b762*16 + a27*28*16] = data_11_array[a27][b762][m762];
        end
    endgenerate
    generate 
        localparam integer b763 = 7;
        for (m763 = 0; m763 < 16; m763 = m763 + 1) 
        begin: inbit763
            assign data_11[m763 + b763*16 + a27*28*16] = data_11_array[a27][b763][m763];
        end
    endgenerate
    generate 
        localparam integer b764 = 8;
        for (m764 = 0; m764 < 16; m764 = m764 + 1) 
        begin: inbit764
            assign data_11[m764 + b764*16 + a27*28*16] = data_11_array[a27][b764][m764];
        end
    endgenerate
    generate 
        localparam integer b765 = 9;
        for (m765 = 0; m765 < 16; m765 = m765 + 1) 
        begin: inbit765
            assign data_11[m765 + b765*16 + a27*28*16] = data_11_array[a27][b765][m765];
        end
    endgenerate
    generate 
        localparam integer b766 = 10;
        for (m766 = 0; m766 < 16; m766 = m766 + 1) 
        begin: inbit766
            assign data_11[m766 + b766*16 + a27*28*16] = data_11_array[a27][b766][m766];
        end
    endgenerate
    generate 
        localparam integer b767 = 11;
        for (m767 = 0; m767 < 16; m767 = m767 + 1) 
        begin: inbit767
            assign data_11[m767 + b767*16 + a27*28*16] = data_11_array[a27][b767][m767];
        end
    endgenerate
    generate 
        localparam integer b768 = 12;
        for (m768 = 0; m768 < 16; m768 = m768 + 1) 
        begin: inbit768
            assign data_11[m768 + b768*16 + a27*28*16] = data_11_array[a27][b768][m768];
        end
    endgenerate
    generate 
        localparam integer b769 = 13;
        for (m769 = 0; m769 < 16; m769 = m769 + 1) 
        begin: inbit769
            assign data_11[m769 + b769*16 + a27*28*16] = data_11_array[a27][b769][m769];
        end
    endgenerate
    generate 
        localparam integer b770 = 14;
        for (m770 = 0; m770 < 16; m770 = m770 + 1) 
        begin: inbit770
            assign data_11[m770 + b770*16 + a27*28*16] = data_11_array[a27][b770][m770];
        end
    endgenerate
    generate 
        localparam integer b771 = 15;
        for (m771 = 0; m771 < 16; m771 = m771 + 1) 
        begin: inbit771
            assign data_11[m771 + b771*16 + a27*28*16] = data_11_array[a27][b771][m771];
        end
    endgenerate
    generate 
        localparam integer b772 = 16;
        for (m772 = 0; m772 < 16; m772 = m772 + 1) 
        begin: inbit772
            assign data_11[m772 + b772*16 + a27*28*16] = data_11_array[a27][b772][m772];
        end
    endgenerate
    generate 
        localparam integer b773 = 17;
        for (m773 = 0; m773 < 16; m773 = m773 + 1) 
        begin: inbit773
            assign data_11[m773 + b773*16 + a27*28*16] = data_11_array[a27][b773][m773];
        end
    endgenerate
    generate 
        localparam integer b774 = 18;
        for (m774 = 0; m774 < 16; m774 = m774 + 1) 
        begin: inbit774
            assign data_11[m774 + b774*16 + a27*28*16] = data_11_array[a27][b774][m774];
        end
    endgenerate
    generate 
        localparam integer b775 = 19;
        for (m775 = 0; m775 < 16; m775 = m775 + 1) 
        begin: inbit775
            assign data_11[m775 + b775*16 + a27*28*16] = data_11_array[a27][b775][m775];
        end
    endgenerate
    generate 
        localparam integer b776 = 20;
        for (m776 = 0; m776 < 16; m776 = m776 + 1) 
        begin: inbit776
            assign data_11[m776 + b776*16 + a27*28*16] = data_11_array[a27][b776][m776];
        end
    endgenerate
    generate 
        localparam integer b777 = 21;
        for (m777 = 0; m777 < 16; m777 = m777 + 1) 
        begin: inbit777
            assign data_11[m777 + b777*16 + a27*28*16] = data_11_array[a27][b777][m777];
        end
    endgenerate
    generate 
        localparam integer b778 = 22;
        for (m778 = 0; m778 < 16; m778 = m778 + 1) 
        begin: inbit778
            assign data_11[m778 + b778*16 + a27*28*16] = data_11_array[a27][b778][m778];
        end
    endgenerate
    generate 
        localparam integer b779 = 23;
        for (m779 = 0; m779 < 16; m779 = m779 + 1) 
        begin: inbit779
            assign data_11[m779 + b779*16 + a27*28*16] = data_11_array[a27][b779][m779];
        end
    endgenerate
    generate 
        localparam integer b780 = 24;
        for (m780 = 0; m780 < 16; m780 = m780 + 1) 
        begin: inbit780
            assign data_11[m780 + b780*16 + a27*28*16] = data_11_array[a27][b780][m780];
        end
    endgenerate
    generate 
        localparam integer b781 = 25;
        for (m781 = 0; m781 < 16; m781 = m781 + 1) 
        begin: inbit781
            assign data_11[m781 + b781*16 + a27*28*16] = data_11_array[a27][b781][m781];
        end
    endgenerate
    generate 
        localparam integer b782 = 26;
        for (m782 = 0; m782 < 16; m782 = m782 + 1) 
        begin: inbit782
            assign data_11[m782 + b782*16 + a27*28*16] = data_11_array[a27][b782][m782];
        end
    endgenerate
    generate 
        localparam integer b783 = 27;
        for (m783 = 0; m783 < 16; m783 = m783 + 1) 
        begin: inbit783
            assign data_11[m783 + b783*16 + a27*28*16] = data_11_array[a27][b783][m783];
        end
    endgenerate
  
  ////ROW 0
  generate
    localparam integer j0 = 0;
    for (i0 = 0; i0 < 24; i0 = i0 + 1)
    begin: addbit0
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j0+0][i0+0]), .Out(multi0[0][i0]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j0+0][i0+1]), .Out(multi0[1][i0]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j0+0][i0+2]), .Out(multi0[2][i0]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j0+0][i0+3]), .Out(multi0[3][i0]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j0+0][i0+4]), .Out(multi0[4][i0]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j0+1][i0+0]), .Out(multi0[5][i0]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j0+1][i0+1]), .Out(multi0[6][i0]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j0+1][i0+2]), .Out(multi0[7][i0]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j0+1][i0+3]), .Out(multi0[8][i0]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j0+1][i0+4]), .Out(multi0[9][i0]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j0+2][i0+0]), .Out(multi0[10][i0]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j0+2][i0+1]), .Out(multi0[11][i0]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j0+2][i0+2]), .Out(multi0[12][i0]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j0+2][i0+3]), .Out(multi0[13][i0]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j0+2][i0+4]), .Out(multi0[14][i0]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j0+3][i0+0]), .Out(multi0[15][i0]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j0+3][i0+1]), .Out(multi0[16][i0]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j0+3][i0+2]), .Out(multi0[17][i0]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j0+3][i0+3]), .Out(multi0[18][i0]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j0+3][i0+4]), .Out(multi0[19][i0]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j0+4][i0+0]), .Out(multi0[20][i0]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j0+4][i0+1]), .Out(multi0[21][i0]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j0+4][i0+2]), .Out(multi0[22][i0]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j0+4][i0+3]), .Out(multi0[23][i0]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j0+4][i0+4]), .Out(multi0[24][i0]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi0[0][i0]), .B(multi0[1][i0]), .Out(sum0[0][i0]));
      FP16_Add stage026(.A(multi0[2][i0]), .B(multi0[3][i0]), .Out(sum0[1][i0]));
      FP16_Add stage027(.A(multi0[4][i0]), .B(multi0[5][i0]), .Out(sum0[2][i0]));
      FP16_Add stage028(.A(multi0[6][i0]), .B(multi0[7][i0]), .Out(sum0[3][i0]));
      FP16_Add stage029(.A(multi0[8][i0]), .B(multi0[9][i0]), .Out(sum0[4][i0]));
      FP16_Add stage030(.A(multi0[10][i0]), .B(multi0[11][i0]), .Out(sum0[5][i0]));
      FP16_Add stage031(.A(multi0[12][i0]), .B(multi0[13][i0]), .Out(sum0[6][i0]));
      FP16_Add stage032(.A(multi0[14][i0]), .B(multi0[15][i0]), .Out(sum0[7][i0]));
      FP16_Add stage033(.A(multi0[16][i0]), .B(multi0[17][i0]), .Out(sum0[8][i0]));
      FP16_Add stage034(.A(multi0[18][i0]), .B(multi0[19][i0]), .Out(sum0[9][i0]));
      FP16_Add stage035(.A(multi0[20][i0]), .B(multi0[21][i0]), .Out(sum0[10][i0]));
      FP16_Add stage036(.A(multi0[22][i0]), .B(multi0[23][i0]), .Out(sum0[11][i0]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum0[0][i0]), .B(sum0[1][i0]), .Out(sum0[12][i0]));
      FP16_Add stage038(.A(sum0[2][i0]), .B(sum0[3][i0]), .Out(sum0[13][i0]));
      FP16_Add stage039(.A(sum0[4][i0]), .B(sum0[5][i0]), .Out(sum0[14][i0]));
      FP16_Add stage040(.A(sum0[6][i0]), .B(sum0[7][i0]), .Out(sum0[15][i0]));
      FP16_Add stage041(.A(sum0[8][i0]), .B(sum0[9][i0]), .Out(sum0[16][i0]));
      FP16_Add stage042(.A(sum0[10][i0]), .B(sum0[11][i0]), .Out(sum0[17][i0]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum0[12][i0]), .B(sum0[13][i0]), .Out(sum0[18][i0]));
      FP16_Add stage044(.A(sum0[14][i0]), .B(sum0[15][i0]), .Out(sum0[19][i0]));
      FP16_Add stage045(.A(sum0[16][i0]), .B(sum0[17][i0]), .Out(sum0[20][i0]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum0[18][i0]), .B(sum0[19][i0]), .Out(sum0[21][i0]));
      FP16_Add stage047(.A(sum0[20][i0]), .B(multi0[24][i0]), .Out(sum0[22][i0]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum0[21][i0]), .B(sum0[22][i0]), .Out(sum0[23][i0]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum0[23][i0]), .B(feature2Bias), .Out(data_11_array[j0][i0]));
    end
  endgenerate
  
  ////ROW 1
  generate
    localparam integer j1 = 1;
    for (i1 = 0; i1 < 24; i1 = i1 + 1)
    begin: addbit1
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j1+0][i1+0]), .Out(multi1[0][i1]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j1+0][i1+1]), .Out(multi1[1][i1]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j1+0][i1+2]), .Out(multi1[2][i1]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j1+0][i1+3]), .Out(multi1[3][i1]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j1+0][i1+4]), .Out(multi1[4][i1]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j1+1][i1+0]), .Out(multi1[5][i1]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j1+1][i1+1]), .Out(multi1[6][i1]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j1+1][i1+2]), .Out(multi1[7][i1]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j1+1][i1+3]), .Out(multi1[8][i1]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j1+1][i1+4]), .Out(multi1[9][i1]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j1+2][i1+0]), .Out(multi1[10][i1]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j1+2][i1+1]), .Out(multi1[11][i1]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j1+2][i1+2]), .Out(multi1[12][i1]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j1+2][i1+3]), .Out(multi1[13][i1]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j1+2][i1+4]), .Out(multi1[14][i1]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j1+3][i1+0]), .Out(multi1[15][i1]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j1+3][i1+1]), .Out(multi1[16][i1]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j1+3][i1+2]), .Out(multi1[17][i1]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j1+3][i1+3]), .Out(multi1[18][i1]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j1+3][i1+4]), .Out(multi1[19][i1]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j1+4][i1+0]), .Out(multi1[20][i1]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j1+4][i1+1]), .Out(multi1[21][i1]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j1+4][i1+2]), .Out(multi1[22][i1]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j1+4][i1+3]), .Out(multi1[23][i1]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j1+4][i1+4]), .Out(multi1[24][i1]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi1[0][i1]), .B(multi1[1][i1]), .Out(sum1[0][i1]));
      FP16_Add stage026(.A(multi1[2][i1]), .B(multi1[3][i1]), .Out(sum1[1][i1]));
      FP16_Add stage027(.A(multi1[4][i1]), .B(multi1[5][i1]), .Out(sum1[2][i1]));
      FP16_Add stage028(.A(multi1[6][i1]), .B(multi1[7][i1]), .Out(sum1[3][i1]));
      FP16_Add stage029(.A(multi1[8][i1]), .B(multi1[9][i1]), .Out(sum1[4][i1]));
      FP16_Add stage030(.A(multi1[10][i1]), .B(multi1[11][i1]), .Out(sum1[5][i1]));
      FP16_Add stage031(.A(multi1[12][i1]), .B(multi1[13][i1]), .Out(sum1[6][i1]));
      FP16_Add stage032(.A(multi1[14][i1]), .B(multi1[15][i1]), .Out(sum1[7][i1]));
      FP16_Add stage033(.A(multi1[16][i1]), .B(multi1[17][i1]), .Out(sum1[8][i1]));
      FP16_Add stage034(.A(multi1[18][i1]), .B(multi1[19][i1]), .Out(sum1[9][i1]));
      FP16_Add stage035(.A(multi1[20][i1]), .B(multi1[21][i1]), .Out(sum1[10][i1]));
      FP16_Add stage036(.A(multi1[22][i1]), .B(multi1[23][i1]), .Out(sum1[11][i1]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum1[0][i1]), .B(sum1[1][i1]), .Out(sum1[12][i1]));
      FP16_Add stage038(.A(sum1[2][i1]), .B(sum1[3][i1]), .Out(sum1[13][i1]));
      FP16_Add stage039(.A(sum1[4][i1]), .B(sum1[5][i1]), .Out(sum1[14][i1]));
      FP16_Add stage040(.A(sum1[6][i1]), .B(sum1[7][i1]), .Out(sum1[15][i1]));
      FP16_Add stage041(.A(sum1[8][i1]), .B(sum1[9][i1]), .Out(sum1[16][i1]));
      FP16_Add stage042(.A(sum1[10][i1]), .B(sum1[11][i1]), .Out(sum1[17][i1]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum1[12][i1]), .B(sum1[13][i1]), .Out(sum1[18][i1]));
      FP16_Add stage044(.A(sum1[14][i1]), .B(sum1[15][i1]), .Out(sum1[19][i1]));
      FP16_Add stage045(.A(sum1[16][i1]), .B(sum1[17][i1]), .Out(sum1[20][i1]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum1[18][i1]), .B(sum1[19][i1]), .Out(sum1[21][i1]));
      FP16_Add stage047(.A(sum1[20][i1]), .B(multi1[24][i1]), .Out(sum1[22][i1]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum1[21][i1]), .B(sum1[22][i1]), .Out(sum1[23][i1]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum1[23][i1]), .B(feature2Bias), .Out(data_11_array[j1][i1]));
    end
  endgenerate
  
  ////ROW 2
  generate
    localparam integer j2 = 2;
    for (i2 = 0; i2 < 24; i2 = i2 + 1)
    begin: addbit2
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j2+0][i2+0]), .Out(multi2[0][i2]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j2+0][i2+1]), .Out(multi2[1][i2]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j2+0][i2+2]), .Out(multi2[2][i2]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j2+0][i2+3]), .Out(multi2[3][i2]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j2+0][i2+4]), .Out(multi2[4][i2]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j2+1][i2+0]), .Out(multi2[5][i2]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j2+1][i2+1]), .Out(multi2[6][i2]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j2+1][i2+2]), .Out(multi2[7][i2]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j2+1][i2+3]), .Out(multi2[8][i2]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j2+1][i2+4]), .Out(multi2[9][i2]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j2+2][i2+0]), .Out(multi2[10][i2]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j2+2][i2+1]), .Out(multi2[11][i2]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j2+2][i2+2]), .Out(multi2[12][i2]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j2+2][i2+3]), .Out(multi2[13][i2]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j2+2][i2+4]), .Out(multi2[14][i2]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j2+3][i2+0]), .Out(multi2[15][i2]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j2+3][i2+1]), .Out(multi2[16][i2]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j2+3][i2+2]), .Out(multi2[17][i2]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j2+3][i2+3]), .Out(multi2[18][i2]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j2+3][i2+4]), .Out(multi2[19][i2]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j2+4][i2+0]), .Out(multi2[20][i2]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j2+4][i2+1]), .Out(multi2[21][i2]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j2+4][i2+2]), .Out(multi2[22][i2]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j2+4][i2+3]), .Out(multi2[23][i2]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j2+4][i2+4]), .Out(multi2[24][i2]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi2[0][i2]), .B(multi2[1][i2]), .Out(sum2[0][i2]));
      FP16_Add stage026(.A(multi2[2][i2]), .B(multi2[3][i2]), .Out(sum2[1][i2]));
      FP16_Add stage027(.A(multi2[4][i2]), .B(multi2[5][i2]), .Out(sum2[2][i2]));
      FP16_Add stage028(.A(multi2[6][i2]), .B(multi2[7][i2]), .Out(sum2[3][i2]));
      FP16_Add stage029(.A(multi2[8][i2]), .B(multi2[9][i2]), .Out(sum2[4][i2]));
      FP16_Add stage030(.A(multi2[10][i2]), .B(multi2[11][i2]), .Out(sum2[5][i2]));
      FP16_Add stage031(.A(multi2[12][i2]), .B(multi2[13][i2]), .Out(sum2[6][i2]));
      FP16_Add stage032(.A(multi2[14][i2]), .B(multi2[15][i2]), .Out(sum2[7][i2]));
      FP16_Add stage033(.A(multi2[16][i2]), .B(multi2[17][i2]), .Out(sum2[8][i2]));
      FP16_Add stage034(.A(multi2[18][i2]), .B(multi2[19][i2]), .Out(sum2[9][i2]));
      FP16_Add stage035(.A(multi2[20][i2]), .B(multi2[21][i2]), .Out(sum2[10][i2]));
      FP16_Add stage036(.A(multi2[22][i2]), .B(multi2[23][i2]), .Out(sum2[11][i2]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum2[0][i2]), .B(sum2[1][i2]), .Out(sum2[12][i2]));
      FP16_Add stage038(.A(sum2[2][i2]), .B(sum2[3][i2]), .Out(sum2[13][i2]));
      FP16_Add stage039(.A(sum2[4][i2]), .B(sum2[5][i2]), .Out(sum2[14][i2]));
      FP16_Add stage040(.A(sum2[6][i2]), .B(sum2[7][i2]), .Out(sum2[15][i2]));
      FP16_Add stage041(.A(sum2[8][i2]), .B(sum2[9][i2]), .Out(sum2[16][i2]));
      FP16_Add stage042(.A(sum2[10][i2]), .B(sum2[11][i2]), .Out(sum2[17][i2]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum2[12][i2]), .B(sum2[13][i2]), .Out(sum2[18][i2]));
      FP16_Add stage044(.A(sum2[14][i2]), .B(sum2[15][i2]), .Out(sum2[19][i2]));
      FP16_Add stage045(.A(sum2[16][i2]), .B(sum2[17][i2]), .Out(sum2[20][i2]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum2[18][i2]), .B(sum2[19][i2]), .Out(sum2[21][i2]));
      FP16_Add stage047(.A(sum2[20][i2]), .B(multi2[24][i2]), .Out(sum2[22][i2]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum2[21][i2]), .B(sum2[22][i2]), .Out(sum2[23][i2]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum2[23][i2]), .B(feature2Bias), .Out(data_11_array[j2][i2]));
    end
  endgenerate
  
  ////ROW 3
  generate
    localparam integer j3 = 3;
    for (i3 = 0; i3 < 24; i3 = i3 + 1)
    begin: addbit3
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j3+0][i3+0]), .Out(multi3[0][i3]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j3+0][i3+1]), .Out(multi3[1][i3]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j3+0][i3+2]), .Out(multi3[2][i3]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j3+0][i3+3]), .Out(multi3[3][i3]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j3+0][i3+4]), .Out(multi3[4][i3]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j3+1][i3+0]), .Out(multi3[5][i3]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j3+1][i3+1]), .Out(multi3[6][i3]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j3+1][i3+2]), .Out(multi3[7][i3]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j3+1][i3+3]), .Out(multi3[8][i3]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j3+1][i3+4]), .Out(multi3[9][i3]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j3+2][i3+0]), .Out(multi3[10][i3]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j3+2][i3+1]), .Out(multi3[11][i3]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j3+2][i3+2]), .Out(multi3[12][i3]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j3+2][i3+3]), .Out(multi3[13][i3]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j3+2][i3+4]), .Out(multi3[14][i3]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j3+3][i3+0]), .Out(multi3[15][i3]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j3+3][i3+1]), .Out(multi3[16][i3]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j3+3][i3+2]), .Out(multi3[17][i3]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j3+3][i3+3]), .Out(multi3[18][i3]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j3+3][i3+4]), .Out(multi3[19][i3]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j3+4][i3+0]), .Out(multi3[20][i3]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j3+4][i3+1]), .Out(multi3[21][i3]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j3+4][i3+2]), .Out(multi3[22][i3]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j3+4][i3+3]), .Out(multi3[23][i3]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j3+4][i3+4]), .Out(multi3[24][i3]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi3[0][i3]), .B(multi3[1][i3]), .Out(sum3[0][i3]));
      FP16_Add stage026(.A(multi3[2][i3]), .B(multi3[3][i3]), .Out(sum3[1][i3]));
      FP16_Add stage027(.A(multi3[4][i3]), .B(multi3[5][i3]), .Out(sum3[2][i3]));
      FP16_Add stage028(.A(multi3[6][i3]), .B(multi3[7][i3]), .Out(sum3[3][i3]));
      FP16_Add stage029(.A(multi3[8][i3]), .B(multi3[9][i3]), .Out(sum3[4][i3]));
      FP16_Add stage030(.A(multi3[10][i3]), .B(multi3[11][i3]), .Out(sum3[5][i3]));
      FP16_Add stage031(.A(multi3[12][i3]), .B(multi3[13][i3]), .Out(sum3[6][i3]));
      FP16_Add stage032(.A(multi3[14][i3]), .B(multi3[15][i3]), .Out(sum3[7][i3]));
      FP16_Add stage033(.A(multi3[16][i3]), .B(multi3[17][i3]), .Out(sum3[8][i3]));
      FP16_Add stage034(.A(multi3[18][i3]), .B(multi3[19][i3]), .Out(sum3[9][i3]));
      FP16_Add stage035(.A(multi3[20][i3]), .B(multi3[21][i3]), .Out(sum3[10][i3]));
      FP16_Add stage036(.A(multi3[22][i3]), .B(multi3[23][i3]), .Out(sum3[11][i3]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum3[0][i3]), .B(sum3[1][i3]), .Out(sum3[12][i3]));
      FP16_Add stage038(.A(sum3[2][i3]), .B(sum3[3][i3]), .Out(sum3[13][i3]));
      FP16_Add stage039(.A(sum3[4][i3]), .B(sum3[5][i3]), .Out(sum3[14][i3]));
      FP16_Add stage040(.A(sum3[6][i3]), .B(sum3[7][i3]), .Out(sum3[15][i3]));
      FP16_Add stage041(.A(sum3[8][i3]), .B(sum3[9][i3]), .Out(sum3[16][i3]));
      FP16_Add stage042(.A(sum3[10][i3]), .B(sum3[11][i3]), .Out(sum3[17][i3]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum3[12][i3]), .B(sum3[13][i3]), .Out(sum3[18][i3]));
      FP16_Add stage044(.A(sum3[14][i3]), .B(sum3[15][i3]), .Out(sum3[19][i3]));
      FP16_Add stage045(.A(sum3[16][i3]), .B(sum3[17][i3]), .Out(sum3[20][i3]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum3[18][i3]), .B(sum3[19][i3]), .Out(sum3[21][i3]));
      FP16_Add stage047(.A(sum3[20][i3]), .B(multi3[24][i3]), .Out(sum3[22][i3]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum3[21][i3]), .B(sum3[22][i3]), .Out(sum3[23][i3]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum3[23][i3]), .B(feature2Bias), .Out(data_11_array[j3][i3]));
    end
  endgenerate
  
  ////ROW 4
  generate
    localparam integer j4 = 4;
    for (i4 = 0; i4 < 24; i4 = i4 + 1)
    begin: addbit4
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j4+0][i4+0]), .Out(multi4[0][i4]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j4+0][i4+1]), .Out(multi4[1][i4]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j4+0][i4+2]), .Out(multi4[2][i4]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j4+0][i4+3]), .Out(multi4[3][i4]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j4+0][i4+4]), .Out(multi4[4][i4]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j4+1][i4+0]), .Out(multi4[5][i4]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j4+1][i4+1]), .Out(multi4[6][i4]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j4+1][i4+2]), .Out(multi4[7][i4]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j4+1][i4+3]), .Out(multi4[8][i4]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j4+1][i4+4]), .Out(multi4[9][i4]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j4+2][i4+0]), .Out(multi4[10][i4]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j4+2][i4+1]), .Out(multi4[11][i4]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j4+2][i4+2]), .Out(multi4[12][i4]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j4+2][i4+3]), .Out(multi4[13][i4]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j4+2][i4+4]), .Out(multi4[14][i4]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j4+3][i4+0]), .Out(multi4[15][i4]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j4+3][i4+1]), .Out(multi4[16][i4]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j4+3][i4+2]), .Out(multi4[17][i4]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j4+3][i4+3]), .Out(multi4[18][i4]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j4+3][i4+4]), .Out(multi4[19][i4]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j4+4][i4+0]), .Out(multi4[20][i4]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j4+4][i4+1]), .Out(multi4[21][i4]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j4+4][i4+2]), .Out(multi4[22][i4]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j4+4][i4+3]), .Out(multi4[23][i4]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j4+4][i4+4]), .Out(multi4[24][i4]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi4[0][i4]), .B(multi4[1][i4]), .Out(sum4[0][i4]));
      FP16_Add stage026(.A(multi4[2][i4]), .B(multi4[3][i4]), .Out(sum4[1][i4]));
      FP16_Add stage027(.A(multi4[4][i4]), .B(multi4[5][i4]), .Out(sum4[2][i4]));
      FP16_Add stage028(.A(multi4[6][i4]), .B(multi4[7][i4]), .Out(sum4[3][i4]));
      FP16_Add stage029(.A(multi4[8][i4]), .B(multi4[9][i4]), .Out(sum4[4][i4]));
      FP16_Add stage030(.A(multi4[10][i4]), .B(multi4[11][i4]), .Out(sum4[5][i4]));
      FP16_Add stage031(.A(multi4[12][i4]), .B(multi4[13][i4]), .Out(sum4[6][i4]));
      FP16_Add stage032(.A(multi4[14][i4]), .B(multi4[15][i4]), .Out(sum4[7][i4]));
      FP16_Add stage033(.A(multi4[16][i4]), .B(multi4[17][i4]), .Out(sum4[8][i4]));
      FP16_Add stage034(.A(multi4[18][i4]), .B(multi4[19][i4]), .Out(sum4[9][i4]));
      FP16_Add stage035(.A(multi4[20][i4]), .B(multi4[21][i4]), .Out(sum4[10][i4]));
      FP16_Add stage036(.A(multi4[22][i4]), .B(multi4[23][i4]), .Out(sum4[11][i4]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum4[0][i4]), .B(sum4[1][i4]), .Out(sum4[12][i4]));
      FP16_Add stage038(.A(sum4[2][i4]), .B(sum4[3][i4]), .Out(sum4[13][i4]));
      FP16_Add stage039(.A(sum4[4][i4]), .B(sum4[5][i4]), .Out(sum4[14][i4]));
      FP16_Add stage040(.A(sum4[6][i4]), .B(sum4[7][i4]), .Out(sum4[15][i4]));
      FP16_Add stage041(.A(sum4[8][i4]), .B(sum4[9][i4]), .Out(sum4[16][i4]));
      FP16_Add stage042(.A(sum4[10][i4]), .B(sum4[11][i4]), .Out(sum4[17][i4]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum4[12][i4]), .B(sum4[13][i4]), .Out(sum4[18][i4]));
      FP16_Add stage044(.A(sum4[14][i4]), .B(sum4[15][i4]), .Out(sum4[19][i4]));
      FP16_Add stage045(.A(sum4[16][i4]), .B(sum4[17][i4]), .Out(sum4[20][i4]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum4[18][i4]), .B(sum4[19][i4]), .Out(sum4[21][i4]));
      FP16_Add stage047(.A(sum4[20][i4]), .B(multi4[24][i4]), .Out(sum4[22][i4]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum4[21][i4]), .B(sum4[22][i4]), .Out(sum4[23][i4]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum4[23][i4]), .B(feature2Bias), .Out(data_11_array[j4][i4]));
    end
  endgenerate
  
  ////ROW 5
  generate
    localparam integer j5 = 5;
    for (i5 = 0; i5 < 24; i5 = i5 + 1)
    begin: addbit5
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j5+0][i5+0]), .Out(multi5[0][i5]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j5+0][i5+1]), .Out(multi5[1][i5]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j5+0][i5+2]), .Out(multi5[2][i5]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j5+0][i5+3]), .Out(multi5[3][i5]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j5+0][i5+4]), .Out(multi5[4][i5]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j5+1][i5+0]), .Out(multi5[5][i5]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j5+1][i5+1]), .Out(multi5[6][i5]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j5+1][i5+2]), .Out(multi5[7][i5]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j5+1][i5+3]), .Out(multi5[8][i5]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j5+1][i5+4]), .Out(multi5[9][i5]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j5+2][i5+0]), .Out(multi5[10][i5]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j5+2][i5+1]), .Out(multi5[11][i5]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j5+2][i5+2]), .Out(multi5[12][i5]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j5+2][i5+3]), .Out(multi5[13][i5]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j5+2][i5+4]), .Out(multi5[14][i5]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j5+3][i5+0]), .Out(multi5[15][i5]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j5+3][i5+1]), .Out(multi5[16][i5]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j5+3][i5+2]), .Out(multi5[17][i5]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j5+3][i5+3]), .Out(multi5[18][i5]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j5+3][i5+4]), .Out(multi5[19][i5]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j5+4][i5+0]), .Out(multi5[20][i5]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j5+4][i5+1]), .Out(multi5[21][i5]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j5+4][i5+2]), .Out(multi5[22][i5]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j5+4][i5+3]), .Out(multi5[23][i5]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j5+4][i5+4]), .Out(multi5[24][i5]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi5[0][i5]), .B(multi5[1][i5]), .Out(sum5[0][i5]));
      FP16_Add stage026(.A(multi5[2][i5]), .B(multi5[3][i5]), .Out(sum5[1][i5]));
      FP16_Add stage027(.A(multi5[4][i5]), .B(multi5[5][i5]), .Out(sum5[2][i5]));
      FP16_Add stage028(.A(multi5[6][i5]), .B(multi5[7][i5]), .Out(sum5[3][i5]));
      FP16_Add stage029(.A(multi5[8][i5]), .B(multi5[9][i5]), .Out(sum5[4][i5]));
      FP16_Add stage030(.A(multi5[10][i5]), .B(multi5[11][i5]), .Out(sum5[5][i5]));
      FP16_Add stage031(.A(multi5[12][i5]), .B(multi5[13][i5]), .Out(sum5[6][i5]));
      FP16_Add stage032(.A(multi5[14][i5]), .B(multi5[15][i5]), .Out(sum5[7][i5]));
      FP16_Add stage033(.A(multi5[16][i5]), .B(multi5[17][i5]), .Out(sum5[8][i5]));
      FP16_Add stage034(.A(multi5[18][i5]), .B(multi5[19][i5]), .Out(sum5[9][i5]));
      FP16_Add stage035(.A(multi5[20][i5]), .B(multi5[21][i5]), .Out(sum5[10][i5]));
      FP16_Add stage036(.A(multi5[22][i5]), .B(multi5[23][i5]), .Out(sum5[11][i5]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum5[0][i5]), .B(sum5[1][i5]), .Out(sum5[12][i5]));
      FP16_Add stage038(.A(sum5[2][i5]), .B(sum5[3][i5]), .Out(sum5[13][i5]));
      FP16_Add stage039(.A(sum5[4][i5]), .B(sum5[5][i5]), .Out(sum5[14][i5]));
      FP16_Add stage040(.A(sum5[6][i5]), .B(sum5[7][i5]), .Out(sum5[15][i5]));
      FP16_Add stage041(.A(sum5[8][i5]), .B(sum5[9][i5]), .Out(sum5[16][i5]));
      FP16_Add stage042(.A(sum5[10][i5]), .B(sum5[11][i5]), .Out(sum5[17][i5]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum5[12][i5]), .B(sum5[13][i5]), .Out(sum5[18][i5]));
      FP16_Add stage044(.A(sum5[14][i5]), .B(sum5[15][i5]), .Out(sum5[19][i5]));
      FP16_Add stage045(.A(sum5[16][i5]), .B(sum5[17][i5]), .Out(sum5[20][i5]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum5[18][i5]), .B(sum5[19][i5]), .Out(sum5[21][i5]));
      FP16_Add stage047(.A(sum5[20][i5]), .B(multi5[24][i5]), .Out(sum5[22][i5]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum5[21][i5]), .B(sum5[22][i5]), .Out(sum5[23][i5]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum5[23][i5]), .B(feature2Bias), .Out(data_11_array[j5][i5]));
    end
  endgenerate
  
  ////ROW 6
  generate
    localparam integer j6 = 6;
    for (i6 = 0; i6 < 24; i6 = i6 + 1)
    begin: addbit6
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j6+0][i6+0]), .Out(multi6[0][i6]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j6+0][i6+1]), .Out(multi6[1][i6]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j6+0][i6+2]), .Out(multi6[2][i6]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j6+0][i6+3]), .Out(multi6[3][i6]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j6+0][i6+4]), .Out(multi6[4][i6]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j6+1][i6+0]), .Out(multi6[5][i6]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j6+1][i6+1]), .Out(multi6[6][i6]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j6+1][i6+2]), .Out(multi6[7][i6]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j6+1][i6+3]), .Out(multi6[8][i6]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j6+1][i6+4]), .Out(multi6[9][i6]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j6+2][i6+0]), .Out(multi6[10][i6]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j6+2][i6+1]), .Out(multi6[11][i6]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j6+2][i6+2]), .Out(multi6[12][i6]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j6+2][i6+3]), .Out(multi6[13][i6]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j6+2][i6+4]), .Out(multi6[14][i6]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j6+3][i6+0]), .Out(multi6[15][i6]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j6+3][i6+1]), .Out(multi6[16][i6]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j6+3][i6+2]), .Out(multi6[17][i6]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j6+3][i6+3]), .Out(multi6[18][i6]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j6+3][i6+4]), .Out(multi6[19][i6]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j6+4][i6+0]), .Out(multi6[20][i6]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j6+4][i6+1]), .Out(multi6[21][i6]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j6+4][i6+2]), .Out(multi6[22][i6]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j6+4][i6+3]), .Out(multi6[23][i6]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j6+4][i6+4]), .Out(multi6[24][i6]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi6[0][i6]), .B(multi6[1][i6]), .Out(sum6[0][i6]));
      FP16_Add stage026(.A(multi6[2][i6]), .B(multi6[3][i6]), .Out(sum6[1][i6]));
      FP16_Add stage027(.A(multi6[4][i6]), .B(multi6[5][i6]), .Out(sum6[2][i6]));
      FP16_Add stage028(.A(multi6[6][i6]), .B(multi6[7][i6]), .Out(sum6[3][i6]));
      FP16_Add stage029(.A(multi6[8][i6]), .B(multi6[9][i6]), .Out(sum6[4][i6]));
      FP16_Add stage030(.A(multi6[10][i6]), .B(multi6[11][i6]), .Out(sum6[5][i6]));
      FP16_Add stage031(.A(multi6[12][i6]), .B(multi6[13][i6]), .Out(sum6[6][i6]));
      FP16_Add stage032(.A(multi6[14][i6]), .B(multi6[15][i6]), .Out(sum6[7][i6]));
      FP16_Add stage033(.A(multi6[16][i6]), .B(multi6[17][i6]), .Out(sum6[8][i6]));
      FP16_Add stage034(.A(multi6[18][i6]), .B(multi6[19][i6]), .Out(sum6[9][i6]));
      FP16_Add stage035(.A(multi6[20][i6]), .B(multi6[21][i6]), .Out(sum6[10][i6]));
      FP16_Add stage036(.A(multi6[22][i6]), .B(multi6[23][i6]), .Out(sum6[11][i6]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum6[0][i6]), .B(sum6[1][i6]), .Out(sum6[12][i6]));
      FP16_Add stage038(.A(sum6[2][i6]), .B(sum6[3][i6]), .Out(sum6[13][i6]));
      FP16_Add stage039(.A(sum6[4][i6]), .B(sum6[5][i6]), .Out(sum6[14][i6]));
      FP16_Add stage040(.A(sum6[6][i6]), .B(sum6[7][i6]), .Out(sum6[15][i6]));
      FP16_Add stage041(.A(sum6[8][i6]), .B(sum6[9][i6]), .Out(sum6[16][i6]));
      FP16_Add stage042(.A(sum6[10][i6]), .B(sum6[11][i6]), .Out(sum6[17][i6]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum6[12][i6]), .B(sum6[13][i6]), .Out(sum6[18][i6]));
      FP16_Add stage044(.A(sum6[14][i6]), .B(sum6[15][i6]), .Out(sum6[19][i6]));
      FP16_Add stage045(.A(sum6[16][i6]), .B(sum6[17][i6]), .Out(sum6[20][i6]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum6[18][i6]), .B(sum6[19][i6]), .Out(sum6[21][i6]));
      FP16_Add stage047(.A(sum6[20][i6]), .B(multi6[24][i6]), .Out(sum6[22][i6]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum6[21][i6]), .B(sum6[22][i6]), .Out(sum6[23][i6]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum6[23][i6]), .B(feature2Bias), .Out(data_11_array[j6][i6]));
    end
  endgenerate
  
  ////ROW 7
  generate
    localparam integer j7 = 7;
    for (i7 = 0; i7 < 24; i7 = i7 + 1)
    begin: addbit7
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j7+0][i7+0]), .Out(multi7[0][i7]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j7+0][i7+1]), .Out(multi7[1][i7]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j7+0][i7+2]), .Out(multi7[2][i7]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j7+0][i7+3]), .Out(multi7[3][i7]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j7+0][i7+4]), .Out(multi7[4][i7]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j7+1][i7+0]), .Out(multi7[5][i7]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j7+1][i7+1]), .Out(multi7[6][i7]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j7+1][i7+2]), .Out(multi7[7][i7]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j7+1][i7+3]), .Out(multi7[8][i7]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j7+1][i7+4]), .Out(multi7[9][i7]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j7+2][i7+0]), .Out(multi7[10][i7]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j7+2][i7+1]), .Out(multi7[11][i7]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j7+2][i7+2]), .Out(multi7[12][i7]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j7+2][i7+3]), .Out(multi7[13][i7]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j7+2][i7+4]), .Out(multi7[14][i7]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j7+3][i7+0]), .Out(multi7[15][i7]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j7+3][i7+1]), .Out(multi7[16][i7]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j7+3][i7+2]), .Out(multi7[17][i7]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j7+3][i7+3]), .Out(multi7[18][i7]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j7+3][i7+4]), .Out(multi7[19][i7]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j7+4][i7+0]), .Out(multi7[20][i7]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j7+4][i7+1]), .Out(multi7[21][i7]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j7+4][i7+2]), .Out(multi7[22][i7]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j7+4][i7+3]), .Out(multi7[23][i7]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j7+4][i7+4]), .Out(multi7[24][i7]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi7[0][i7]), .B(multi7[1][i7]), .Out(sum7[0][i7]));
      FP16_Add stage026(.A(multi7[2][i7]), .B(multi7[3][i7]), .Out(sum7[1][i7]));
      FP16_Add stage027(.A(multi7[4][i7]), .B(multi7[5][i7]), .Out(sum7[2][i7]));
      FP16_Add stage028(.A(multi7[6][i7]), .B(multi7[7][i7]), .Out(sum7[3][i7]));
      FP16_Add stage029(.A(multi7[8][i7]), .B(multi7[9][i7]), .Out(sum7[4][i7]));
      FP16_Add stage030(.A(multi7[10][i7]), .B(multi7[11][i7]), .Out(sum7[5][i7]));
      FP16_Add stage031(.A(multi7[12][i7]), .B(multi7[13][i7]), .Out(sum7[6][i7]));
      FP16_Add stage032(.A(multi7[14][i7]), .B(multi7[15][i7]), .Out(sum7[7][i7]));
      FP16_Add stage033(.A(multi7[16][i7]), .B(multi7[17][i7]), .Out(sum7[8][i7]));
      FP16_Add stage034(.A(multi7[18][i7]), .B(multi7[19][i7]), .Out(sum7[9][i7]));
      FP16_Add stage035(.A(multi7[20][i7]), .B(multi7[21][i7]), .Out(sum7[10][i7]));
      FP16_Add stage036(.A(multi7[22][i7]), .B(multi7[23][i7]), .Out(sum7[11][i7]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum7[0][i7]), .B(sum7[1][i7]), .Out(sum7[12][i7]));
      FP16_Add stage038(.A(sum7[2][i7]), .B(sum7[3][i7]), .Out(sum7[13][i7]));
      FP16_Add stage039(.A(sum7[4][i7]), .B(sum7[5][i7]), .Out(sum7[14][i7]));
      FP16_Add stage040(.A(sum7[6][i7]), .B(sum7[7][i7]), .Out(sum7[15][i7]));
      FP16_Add stage041(.A(sum7[8][i7]), .B(sum7[9][i7]), .Out(sum7[16][i7]));
      FP16_Add stage042(.A(sum7[10][i7]), .B(sum7[11][i7]), .Out(sum7[17][i7]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum7[12][i7]), .B(sum7[13][i7]), .Out(sum7[18][i7]));
      FP16_Add stage044(.A(sum7[14][i7]), .B(sum7[15][i7]), .Out(sum7[19][i7]));
      FP16_Add stage045(.A(sum7[16][i7]), .B(sum7[17][i7]), .Out(sum7[20][i7]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum7[18][i7]), .B(sum7[19][i7]), .Out(sum7[21][i7]));
      FP16_Add stage047(.A(sum7[20][i7]), .B(multi7[24][i7]), .Out(sum7[22][i7]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum7[21][i7]), .B(sum7[22][i7]), .Out(sum7[23][i7]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum7[23][i7]), .B(feature2Bias), .Out(data_11_array[j7][i7]));
    end
  endgenerate
  
  ////ROW 8
  generate
    localparam integer j8 = 8;
    for (i8 = 0; i8 < 24; i8 = i8 + 1)
    begin: addbit8
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j8+0][i8+0]), .Out(multi8[0][i8]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j8+0][i8+1]), .Out(multi8[1][i8]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j8+0][i8+2]), .Out(multi8[2][i8]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j8+0][i8+3]), .Out(multi8[3][i8]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j8+0][i8+4]), .Out(multi8[4][i8]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j8+1][i8+0]), .Out(multi8[5][i8]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j8+1][i8+1]), .Out(multi8[6][i8]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j8+1][i8+2]), .Out(multi8[7][i8]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j8+1][i8+3]), .Out(multi8[8][i8]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j8+1][i8+4]), .Out(multi8[9][i8]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j8+2][i8+0]), .Out(multi8[10][i8]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j8+2][i8+1]), .Out(multi8[11][i8]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j8+2][i8+2]), .Out(multi8[12][i8]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j8+2][i8+3]), .Out(multi8[13][i8]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j8+2][i8+4]), .Out(multi8[14][i8]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j8+3][i8+0]), .Out(multi8[15][i8]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j8+3][i8+1]), .Out(multi8[16][i8]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j8+3][i8+2]), .Out(multi8[17][i8]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j8+3][i8+3]), .Out(multi8[18][i8]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j8+3][i8+4]), .Out(multi8[19][i8]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j8+4][i8+0]), .Out(multi8[20][i8]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j8+4][i8+1]), .Out(multi8[21][i8]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j8+4][i8+2]), .Out(multi8[22][i8]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j8+4][i8+3]), .Out(multi8[23][i8]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j8+4][i8+4]), .Out(multi8[24][i8]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi8[0][i8]), .B(multi8[1][i8]), .Out(sum8[0][i8]));
      FP16_Add stage026(.A(multi8[2][i8]), .B(multi8[3][i8]), .Out(sum8[1][i8]));
      FP16_Add stage027(.A(multi8[4][i8]), .B(multi8[5][i8]), .Out(sum8[2][i8]));
      FP16_Add stage028(.A(multi8[6][i8]), .B(multi8[7][i8]), .Out(sum8[3][i8]));
      FP16_Add stage029(.A(multi8[8][i8]), .B(multi8[9][i8]), .Out(sum8[4][i8]));
      FP16_Add stage030(.A(multi8[10][i8]), .B(multi8[11][i8]), .Out(sum8[5][i8]));
      FP16_Add stage031(.A(multi8[12][i8]), .B(multi8[13][i8]), .Out(sum8[6][i8]));
      FP16_Add stage032(.A(multi8[14][i8]), .B(multi8[15][i8]), .Out(sum8[7][i8]));
      FP16_Add stage033(.A(multi8[16][i8]), .B(multi8[17][i8]), .Out(sum8[8][i8]));
      FP16_Add stage034(.A(multi8[18][i8]), .B(multi8[19][i8]), .Out(sum8[9][i8]));
      FP16_Add stage035(.A(multi8[20][i8]), .B(multi8[21][i8]), .Out(sum8[10][i8]));
      FP16_Add stage036(.A(multi8[22][i8]), .B(multi8[23][i8]), .Out(sum8[11][i8]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum8[0][i8]), .B(sum8[1][i8]), .Out(sum8[12][i8]));
      FP16_Add stage038(.A(sum8[2][i8]), .B(sum8[3][i8]), .Out(sum8[13][i8]));
      FP16_Add stage039(.A(sum8[4][i8]), .B(sum8[5][i8]), .Out(sum8[14][i8]));
      FP16_Add stage040(.A(sum8[6][i8]), .B(sum8[7][i8]), .Out(sum8[15][i8]));
      FP16_Add stage041(.A(sum8[8][i8]), .B(sum8[9][i8]), .Out(sum8[16][i8]));
      FP16_Add stage042(.A(sum8[10][i8]), .B(sum8[11][i8]), .Out(sum8[17][i8]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum8[12][i8]), .B(sum8[13][i8]), .Out(sum8[18][i8]));
      FP16_Add stage044(.A(sum8[14][i8]), .B(sum8[15][i8]), .Out(sum8[19][i8]));
      FP16_Add stage045(.A(sum8[16][i8]), .B(sum8[17][i8]), .Out(sum8[20][i8]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum8[18][i8]), .B(sum8[19][i8]), .Out(sum8[21][i8]));
      FP16_Add stage047(.A(sum8[20][i8]), .B(multi8[24][i8]), .Out(sum8[22][i8]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum8[21][i8]), .B(sum8[22][i8]), .Out(sum8[23][i8]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum8[23][i8]), .B(feature2Bias), .Out(data_11_array[j8][i8]));
    end
  endgenerate
  
  ////ROW 9
  generate
    localparam integer j9 = 9;
    for (i9 = 0; i9 < 24; i9 = i9 + 1)
    begin: addbit9
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j9+0][i9+0]), .Out(multi9[0][i9]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j9+0][i9+1]), .Out(multi9[1][i9]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j9+0][i9+2]), .Out(multi9[2][i9]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j9+0][i9+3]), .Out(multi9[3][i9]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j9+0][i9+4]), .Out(multi9[4][i9]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j9+1][i9+0]), .Out(multi9[5][i9]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j9+1][i9+1]), .Out(multi9[6][i9]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j9+1][i9+2]), .Out(multi9[7][i9]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j9+1][i9+3]), .Out(multi9[8][i9]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j9+1][i9+4]), .Out(multi9[9][i9]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j9+2][i9+0]), .Out(multi9[10][i9]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j9+2][i9+1]), .Out(multi9[11][i9]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j9+2][i9+2]), .Out(multi9[12][i9]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j9+2][i9+3]), .Out(multi9[13][i9]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j9+2][i9+4]), .Out(multi9[14][i9]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j9+3][i9+0]), .Out(multi9[15][i9]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j9+3][i9+1]), .Out(multi9[16][i9]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j9+3][i9+2]), .Out(multi9[17][i9]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j9+3][i9+3]), .Out(multi9[18][i9]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j9+3][i9+4]), .Out(multi9[19][i9]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j9+4][i9+0]), .Out(multi9[20][i9]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j9+4][i9+1]), .Out(multi9[21][i9]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j9+4][i9+2]), .Out(multi9[22][i9]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j9+4][i9+3]), .Out(multi9[23][i9]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j9+4][i9+4]), .Out(multi9[24][i9]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi9[0][i9]), .B(multi9[1][i9]), .Out(sum9[0][i9]));
      FP16_Add stage026(.A(multi9[2][i9]), .B(multi9[3][i9]), .Out(sum9[1][i9]));
      FP16_Add stage027(.A(multi9[4][i9]), .B(multi9[5][i9]), .Out(sum9[2][i9]));
      FP16_Add stage028(.A(multi9[6][i9]), .B(multi9[7][i9]), .Out(sum9[3][i9]));
      FP16_Add stage029(.A(multi9[8][i9]), .B(multi9[9][i9]), .Out(sum9[4][i9]));
      FP16_Add stage030(.A(multi9[10][i9]), .B(multi9[11][i9]), .Out(sum9[5][i9]));
      FP16_Add stage031(.A(multi9[12][i9]), .B(multi9[13][i9]), .Out(sum9[6][i9]));
      FP16_Add stage032(.A(multi9[14][i9]), .B(multi9[15][i9]), .Out(sum9[7][i9]));
      FP16_Add stage033(.A(multi9[16][i9]), .B(multi9[17][i9]), .Out(sum9[8][i9]));
      FP16_Add stage034(.A(multi9[18][i9]), .B(multi9[19][i9]), .Out(sum9[9][i9]));
      FP16_Add stage035(.A(multi9[20][i9]), .B(multi9[21][i9]), .Out(sum9[10][i9]));
      FP16_Add stage036(.A(multi9[22][i9]), .B(multi9[23][i9]), .Out(sum9[11][i9]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum9[0][i9]), .B(sum9[1][i9]), .Out(sum9[12][i9]));
      FP16_Add stage038(.A(sum9[2][i9]), .B(sum9[3][i9]), .Out(sum9[13][i9]));
      FP16_Add stage039(.A(sum9[4][i9]), .B(sum9[5][i9]), .Out(sum9[14][i9]));
      FP16_Add stage040(.A(sum9[6][i9]), .B(sum9[7][i9]), .Out(sum9[15][i9]));
      FP16_Add stage041(.A(sum9[8][i9]), .B(sum9[9][i9]), .Out(sum9[16][i9]));
      FP16_Add stage042(.A(sum9[10][i9]), .B(sum9[11][i9]), .Out(sum9[17][i9]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum9[12][i9]), .B(sum9[13][i9]), .Out(sum9[18][i9]));
      FP16_Add stage044(.A(sum9[14][i9]), .B(sum9[15][i9]), .Out(sum9[19][i9]));
      FP16_Add stage045(.A(sum9[16][i9]), .B(sum9[17][i9]), .Out(sum9[20][i9]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum9[18][i9]), .B(sum9[19][i9]), .Out(sum9[21][i9]));
      FP16_Add stage047(.A(sum9[20][i9]), .B(multi9[24][i9]), .Out(sum9[22][i9]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum9[21][i9]), .B(sum9[22][i9]), .Out(sum9[23][i9]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum9[23][i9]), .B(feature2Bias), .Out(data_11_array[j9][i9]));
    end
  endgenerate
  
  ////ROW 10
  generate
    localparam integer j10 = 10;
    for (i10 = 0; i10 < 24; i10 = i10 + 1)
    begin: addbit10
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j10+0][i10+0]), .Out(multi10[0][i10]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j10+0][i10+1]), .Out(multi10[1][i10]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j10+0][i10+2]), .Out(multi10[2][i10]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j10+0][i10+3]), .Out(multi10[3][i10]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j10+0][i10+4]), .Out(multi10[4][i10]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j10+1][i10+0]), .Out(multi10[5][i10]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j10+1][i10+1]), .Out(multi10[6][i10]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j10+1][i10+2]), .Out(multi10[7][i10]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j10+1][i10+3]), .Out(multi10[8][i10]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j10+1][i10+4]), .Out(multi10[9][i10]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j10+2][i10+0]), .Out(multi10[10][i10]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j10+2][i10+1]), .Out(multi10[11][i10]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j10+2][i10+2]), .Out(multi10[12][i10]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j10+2][i10+3]), .Out(multi10[13][i10]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j10+2][i10+4]), .Out(multi10[14][i10]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j10+3][i10+0]), .Out(multi10[15][i10]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j10+3][i10+1]), .Out(multi10[16][i10]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j10+3][i10+2]), .Out(multi10[17][i10]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j10+3][i10+3]), .Out(multi10[18][i10]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j10+3][i10+4]), .Out(multi10[19][i10]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j10+4][i10+0]), .Out(multi10[20][i10]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j10+4][i10+1]), .Out(multi10[21][i10]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j10+4][i10+2]), .Out(multi10[22][i10]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j10+4][i10+3]), .Out(multi10[23][i10]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j10+4][i10+4]), .Out(multi10[24][i10]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi10[0][i10]), .B(multi10[1][i10]), .Out(sum10[0][i10]));
      FP16_Add stage026(.A(multi10[2][i10]), .B(multi10[3][i10]), .Out(sum10[1][i10]));
      FP16_Add stage027(.A(multi10[4][i10]), .B(multi10[5][i10]), .Out(sum10[2][i10]));
      FP16_Add stage028(.A(multi10[6][i10]), .B(multi10[7][i10]), .Out(sum10[3][i10]));
      FP16_Add stage029(.A(multi10[8][i10]), .B(multi10[9][i10]), .Out(sum10[4][i10]));
      FP16_Add stage030(.A(multi10[10][i10]), .B(multi10[11][i10]), .Out(sum10[5][i10]));
      FP16_Add stage031(.A(multi10[12][i10]), .B(multi10[13][i10]), .Out(sum10[6][i10]));
      FP16_Add stage032(.A(multi10[14][i10]), .B(multi10[15][i10]), .Out(sum10[7][i10]));
      FP16_Add stage033(.A(multi10[16][i10]), .B(multi10[17][i10]), .Out(sum10[8][i10]));
      FP16_Add stage034(.A(multi10[18][i10]), .B(multi10[19][i10]), .Out(sum10[9][i10]));
      FP16_Add stage035(.A(multi10[20][i10]), .B(multi10[21][i10]), .Out(sum10[10][i10]));
      FP16_Add stage036(.A(multi10[22][i10]), .B(multi10[23][i10]), .Out(sum10[11][i10]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum10[0][i10]), .B(sum10[1][i10]), .Out(sum10[12][i10]));
      FP16_Add stage038(.A(sum10[2][i10]), .B(sum10[3][i10]), .Out(sum10[13][i10]));
      FP16_Add stage039(.A(sum10[4][i10]), .B(sum10[5][i10]), .Out(sum10[14][i10]));
      FP16_Add stage040(.A(sum10[6][i10]), .B(sum10[7][i10]), .Out(sum10[15][i10]));
      FP16_Add stage041(.A(sum10[8][i10]), .B(sum10[9][i10]), .Out(sum10[16][i10]));
      FP16_Add stage042(.A(sum10[10][i10]), .B(sum10[11][i10]), .Out(sum10[17][i10]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum10[12][i10]), .B(sum10[13][i10]), .Out(sum10[18][i10]));
      FP16_Add stage044(.A(sum10[14][i10]), .B(sum10[15][i10]), .Out(sum10[19][i10]));
      FP16_Add stage045(.A(sum10[16][i10]), .B(sum10[17][i10]), .Out(sum10[20][i10]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum10[18][i10]), .B(sum10[19][i10]), .Out(sum10[21][i10]));
      FP16_Add stage047(.A(sum10[20][i10]), .B(multi10[24][i10]), .Out(sum10[22][i10]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum10[21][i10]), .B(sum10[22][i10]), .Out(sum10[23][i10]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum10[23][i10]), .B(feature2Bias), .Out(data_11_array[j10][i10]));
    end
  endgenerate
  
    ////ROW 11
  generate
    localparam integer j11 = 11;
    for (i11 = 0; i11 < 24; i11 = i11 + 1)
    begin: addbit11
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j11+0][i11+0]), .Out(multi11[0][i11]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j11+0][i11+1]), .Out(multi11[1][i11]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j11+0][i11+2]), .Out(multi11[2][i11]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j11+0][i11+3]), .Out(multi11[3][i11]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j11+0][i11+4]), .Out(multi11[4][i11]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j11+1][i11+0]), .Out(multi11[5][i11]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j11+1][i11+1]), .Out(multi11[6][i11]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j11+1][i11+2]), .Out(multi11[7][i11]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j11+1][i11+3]), .Out(multi11[8][i11]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j11+1][i11+4]), .Out(multi11[9][i11]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j11+2][i11+0]), .Out(multi11[10][i11]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j11+2][i11+1]), .Out(multi11[11][i11]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j11+2][i11+2]), .Out(multi11[12][i11]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j11+2][i11+3]), .Out(multi11[13][i11]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j11+2][i11+4]), .Out(multi11[14][i11]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j11+3][i11+0]), .Out(multi11[15][i11]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j11+3][i11+1]), .Out(multi11[16][i11]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j11+3][i11+2]), .Out(multi11[17][i11]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j11+3][i11+3]), .Out(multi11[18][i11]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j11+3][i11+4]), .Out(multi11[19][i11]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j11+4][i11+0]), .Out(multi11[20][i11]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j11+4][i11+1]), .Out(multi11[21][i11]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j11+4][i11+2]), .Out(multi11[22][i11]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j11+4][i11+3]), .Out(multi11[23][i11]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j11+4][i11+4]), .Out(multi11[24][i11]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi11[0][i11]), .B(multi11[1][i11]), .Out(sum11[0][i11]));
      FP16_Add stage026(.A(multi11[2][i11]), .B(multi11[3][i11]), .Out(sum11[1][i11]));
      FP16_Add stage027(.A(multi11[4][i11]), .B(multi11[5][i11]), .Out(sum11[2][i11]));
      FP16_Add stage028(.A(multi11[6][i11]), .B(multi11[7][i11]), .Out(sum11[3][i11]));
      FP16_Add stage029(.A(multi11[8][i11]), .B(multi11[9][i11]), .Out(sum11[4][i11]));
      FP16_Add stage030(.A(multi11[10][i11]), .B(multi11[11][i11]), .Out(sum11[5][i11]));
      FP16_Add stage031(.A(multi11[12][i11]), .B(multi11[13][i11]), .Out(sum11[6][i11]));
      FP16_Add stage032(.A(multi11[14][i11]), .B(multi11[15][i11]), .Out(sum11[7][i11]));
      FP16_Add stage033(.A(multi11[16][i11]), .B(multi11[17][i11]), .Out(sum11[8][i11]));
      FP16_Add stage034(.A(multi11[18][i11]), .B(multi11[19][i11]), .Out(sum11[9][i11]));
      FP16_Add stage035(.A(multi11[20][i11]), .B(multi11[21][i11]), .Out(sum11[10][i11]));
      FP16_Add stage036(.A(multi11[22][i11]), .B(multi11[23][i11]), .Out(sum11[11][i11]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum11[0][i11]), .B(sum11[1][i11]), .Out(sum11[12][i11]));
      FP16_Add stage038(.A(sum11[2][i11]), .B(sum11[3][i11]), .Out(sum11[13][i11]));
      FP16_Add stage039(.A(sum11[4][i11]), .B(sum11[5][i11]), .Out(sum11[14][i11]));
      FP16_Add stage040(.A(sum11[6][i11]), .B(sum11[7][i11]), .Out(sum11[15][i11]));
      FP16_Add stage041(.A(sum11[8][i11]), .B(sum11[9][i11]), .Out(sum11[16][i11]));
      FP16_Add stage042(.A(sum11[10][i11]), .B(sum11[11][i11]), .Out(sum11[17][i11]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum11[12][i11]), .B(sum11[13][i11]), .Out(sum11[18][i11]));
      FP16_Add stage044(.A(sum11[14][i11]), .B(sum11[15][i11]), .Out(sum11[19][i11]));
      FP16_Add stage045(.A(sum11[16][i11]), .B(sum11[17][i11]), .Out(sum11[20][i11]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum11[18][i11]), .B(sum11[19][i11]), .Out(sum11[21][i11]));
      FP16_Add stage047(.A(sum11[20][i11]), .B(multi11[24][i11]), .Out(sum11[22][i11]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum11[21][i11]), .B(sum11[22][i11]), .Out(sum11[23][i11]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum11[23][i11]), .B(feature2Bias), .Out(data_11_array[j11][i11]));
    end
  endgenerate

  ////ROW 12
  generate
    localparam integer j12 = 12;
    for (i12 = 0; i12 < 24; i12 = i12 + 1)
    begin: addbit12
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j12+0][i12+0]), .Out(multi12[0][i12]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j12+0][i12+1]), .Out(multi12[1][i12]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j12+0][i12+2]), .Out(multi12[2][i12]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j12+0][i12+3]), .Out(multi12[3][i12]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j12+0][i12+4]), .Out(multi12[4][i12]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j12+1][i12+0]), .Out(multi12[5][i12]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j12+1][i12+1]), .Out(multi12[6][i12]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j12+1][i12+2]), .Out(multi12[7][i12]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j12+1][i12+3]), .Out(multi12[8][i12]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j12+1][i12+4]), .Out(multi12[9][i12]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j12+2][i12+0]), .Out(multi12[10][i12]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j12+2][i12+1]), .Out(multi12[11][i12]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j12+2][i12+2]), .Out(multi12[12][i12]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j12+2][i12+3]), .Out(multi12[13][i12]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j12+2][i12+4]), .Out(multi12[14][i12]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j12+3][i12+0]), .Out(multi12[15][i12]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j12+3][i12+1]), .Out(multi12[16][i12]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j12+3][i12+2]), .Out(multi12[17][i12]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j12+3][i12+3]), .Out(multi12[18][i12]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j12+3][i12+4]), .Out(multi12[19][i12]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j12+4][i12+0]), .Out(multi12[20][i12]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j12+4][i12+1]), .Out(multi12[21][i12]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j12+4][i12+2]), .Out(multi12[22][i12]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j12+4][i12+3]), .Out(multi12[23][i12]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j12+4][i12+4]), .Out(multi12[24][i12]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi12[0][i12]), .B(multi12[1][i12]), .Out(sum12[0][i12]));
      FP16_Add stage026(.A(multi12[2][i12]), .B(multi12[3][i12]), .Out(sum12[1][i12]));
      FP16_Add stage027(.A(multi12[4][i12]), .B(multi12[5][i12]), .Out(sum12[2][i12]));
      FP16_Add stage028(.A(multi12[6][i12]), .B(multi12[7][i12]), .Out(sum12[3][i12]));
      FP16_Add stage029(.A(multi12[8][i12]), .B(multi12[9][i12]), .Out(sum12[4][i12]));
      FP16_Add stage030(.A(multi12[10][i12]), .B(multi12[11][i12]), .Out(sum12[5][i12]));
      FP16_Add stage031(.A(multi12[12][i12]), .B(multi12[13][i12]), .Out(sum12[6][i12]));
      FP16_Add stage032(.A(multi12[14][i12]), .B(multi12[15][i12]), .Out(sum12[7][i12]));
      FP16_Add stage033(.A(multi12[16][i12]), .B(multi12[17][i12]), .Out(sum12[8][i12]));
      FP16_Add stage034(.A(multi12[18][i12]), .B(multi12[19][i12]), .Out(sum12[9][i12]));
      FP16_Add stage035(.A(multi12[20][i12]), .B(multi12[21][i12]), .Out(sum12[10][i12]));
      FP16_Add stage036(.A(multi12[22][i12]), .B(multi12[23][i12]), .Out(sum12[11][i12]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum12[0][i12]), .B(sum12[1][i12]), .Out(sum12[12][i12]));
      FP16_Add stage038(.A(sum12[2][i12]), .B(sum12[3][i12]), .Out(sum12[13][i12]));
      FP16_Add stage039(.A(sum12[4][i12]), .B(sum12[5][i12]), .Out(sum12[14][i12]));
      FP16_Add stage040(.A(sum12[6][i12]), .B(sum12[7][i12]), .Out(sum12[15][i12]));
      FP16_Add stage041(.A(sum12[8][i12]), .B(sum12[9][i12]), .Out(sum12[16][i12]));
      FP16_Add stage042(.A(sum12[10][i12]), .B(sum12[11][i12]), .Out(sum12[17][i12]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum12[12][i12]), .B(sum12[13][i12]), .Out(sum12[18][i12]));
      FP16_Add stage044(.A(sum12[14][i12]), .B(sum12[15][i12]), .Out(sum12[19][i12]));
      FP16_Add stage045(.A(sum12[16][i12]), .B(sum12[17][i12]), .Out(sum12[20][i12]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum12[18][i12]), .B(sum12[19][i12]), .Out(sum12[21][i12]));
      FP16_Add stage047(.A(sum12[20][i12]), .B(multi12[24][i12]), .Out(sum12[22][i12]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum12[21][i12]), .B(sum12[22][i12]), .Out(sum12[23][i12]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum12[23][i12]), .B(feature2Bias), .Out(data_11_array[j12][i12]));
    end
  endgenerate

  ////ROW 13
  generate
    localparam integer j13 = 13;
    for (i13 = 0; i13 < 24; i13 = i13 + 1)
    begin: addbit13
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j13+0][i13+0]), .Out(multi13[0][i13]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j13+0][i13+1]), .Out(multi13[1][i13]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j13+0][i13+2]), .Out(multi13[2][i13]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j13+0][i13+3]), .Out(multi13[3][i13]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j13+0][i13+4]), .Out(multi13[4][i13]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j13+1][i13+0]), .Out(multi13[5][i13]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j13+1][i13+1]), .Out(multi13[6][i13]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j13+1][i13+2]), .Out(multi13[7][i13]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j13+1][i13+3]), .Out(multi13[8][i13]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j13+1][i13+4]), .Out(multi13[9][i13]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j13+2][i13+0]), .Out(multi13[10][i13]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j13+2][i13+1]), .Out(multi13[11][i13]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j13+2][i13+2]), .Out(multi13[12][i13]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j13+2][i13+3]), .Out(multi13[13][i13]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j13+2][i13+4]), .Out(multi13[14][i13]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j13+3][i13+0]), .Out(multi13[15][i13]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j13+3][i13+1]), .Out(multi13[16][i13]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j13+3][i13+2]), .Out(multi13[17][i13]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j13+3][i13+3]), .Out(multi13[18][i13]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j13+3][i13+4]), .Out(multi13[19][i13]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j13+4][i13+0]), .Out(multi13[20][i13]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j13+4][i13+1]), .Out(multi13[21][i13]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j13+4][i13+2]), .Out(multi13[22][i13]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j13+4][i13+3]), .Out(multi13[23][i13]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j13+4][i13+4]), .Out(multi13[24][i13]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi13[0][i13]), .B(multi13[1][i13]), .Out(sum13[0][i13]));
      FP16_Add stage026(.A(multi13[2][i13]), .B(multi13[3][i13]), .Out(sum13[1][i13]));
      FP16_Add stage027(.A(multi13[4][i13]), .B(multi13[5][i13]), .Out(sum13[2][i13]));
      FP16_Add stage028(.A(multi13[6][i13]), .B(multi13[7][i13]), .Out(sum13[3][i13]));
      FP16_Add stage029(.A(multi13[8][i13]), .B(multi13[9][i13]), .Out(sum13[4][i13]));
      FP16_Add stage030(.A(multi13[10][i13]), .B(multi13[11][i13]), .Out(sum13[5][i13]));
      FP16_Add stage031(.A(multi13[12][i13]), .B(multi13[13][i13]), .Out(sum13[6][i13]));
      FP16_Add stage032(.A(multi13[14][i13]), .B(multi13[15][i13]), .Out(sum13[7][i13]));
      FP16_Add stage033(.A(multi13[16][i13]), .B(multi13[17][i13]), .Out(sum13[8][i13]));
      FP16_Add stage034(.A(multi13[18][i13]), .B(multi13[19][i13]), .Out(sum13[9][i13]));
      FP16_Add stage035(.A(multi13[20][i13]), .B(multi13[21][i13]), .Out(sum13[10][i13]));
      FP16_Add stage036(.A(multi13[22][i13]), .B(multi13[23][i13]), .Out(sum13[11][i13]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum13[0][i13]), .B(sum13[1][i13]), .Out(sum13[12][i13]));
      FP16_Add stage038(.A(sum13[2][i13]), .B(sum13[3][i13]), .Out(sum13[13][i13]));
      FP16_Add stage039(.A(sum13[4][i13]), .B(sum13[5][i13]), .Out(sum13[14][i13]));
      FP16_Add stage040(.A(sum13[6][i13]), .B(sum13[7][i13]), .Out(sum13[15][i13]));
      FP16_Add stage041(.A(sum13[8][i13]), .B(sum13[9][i13]), .Out(sum13[16][i13]));
      FP16_Add stage042(.A(sum13[10][i13]), .B(sum13[11][i13]), .Out(sum13[17][i13]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum13[12][i13]), .B(sum13[13][i13]), .Out(sum13[18][i13]));
      FP16_Add stage044(.A(sum13[14][i13]), .B(sum13[15][i13]), .Out(sum13[19][i13]));
      FP16_Add stage045(.A(sum13[16][i13]), .B(sum13[17][i13]), .Out(sum13[20][i13]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum13[18][i13]), .B(sum13[19][i13]), .Out(sum13[21][i13]));
      FP16_Add stage047(.A(sum13[20][i13]), .B(multi13[24][i13]), .Out(sum13[22][i13]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum13[21][i13]), .B(sum13[22][i13]), .Out(sum13[23][i13]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum13[23][i13]), .B(feature2Bias), .Out(data_11_array[j13][i13]));
    end
  endgenerate

  ////ROW 014
  generate
    localparam integer j14 = 14;
    for (i14 = 0; i14 < 24; i14 = i14 + 1)
    begin: addbit14
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j14+0][i14+0]), .Out(multi14[0][i14]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j14+0][i14+1]), .Out(multi14[1][i14]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j14+0][i14+2]), .Out(multi14[2][i14]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j14+0][i14+3]), .Out(multi14[3][i14]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j14+0][i14+4]), .Out(multi14[4][i14]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j14+1][i14+0]), .Out(multi14[5][i14]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j14+1][i14+1]), .Out(multi14[6][i14]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j14+1][i14+2]), .Out(multi14[7][i14]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j14+1][i14+3]), .Out(multi14[8][i14]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j14+1][i14+4]), .Out(multi14[9][i14]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j14+2][i14+0]), .Out(multi14[10][i14]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j14+2][i14+1]), .Out(multi14[11][i14]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j14+2][i14+2]), .Out(multi14[12][i14]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j14+2][i14+3]), .Out(multi14[13][i14]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j14+2][i14+4]), .Out(multi14[14][i14]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j14+3][i14+0]), .Out(multi14[15][i14]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j14+3][i14+1]), .Out(multi14[16][i14]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j14+3][i14+2]), .Out(multi14[17][i14]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j14+3][i14+3]), .Out(multi14[18][i14]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j14+3][i14+4]), .Out(multi14[19][i14]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j14+4][i14+0]), .Out(multi14[20][i14]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j14+4][i14+1]), .Out(multi14[21][i14]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j14+4][i14+2]), .Out(multi14[22][i14]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j14+4][i14+3]), .Out(multi14[23][i14]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j14+4][i14+4]), .Out(multi14[24][i14]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi14[0][i14]), .B(multi14[1][i14]), .Out(sum14[0][i14]));
      FP16_Add stage026(.A(multi14[2][i14]), .B(multi14[3][i14]), .Out(sum14[1][i14]));
      FP16_Add stage027(.A(multi14[4][i14]), .B(multi14[5][i14]), .Out(sum14[2][i14]));
      FP16_Add stage028(.A(multi14[6][i14]), .B(multi14[7][i14]), .Out(sum14[3][i14]));
      FP16_Add stage029(.A(multi14[8][i14]), .B(multi14[9][i14]), .Out(sum14[4][i14]));
      FP16_Add stage030(.A(multi14[10][i14]), .B(multi14[11][i14]), .Out(sum14[5][i14]));
      FP16_Add stage031(.A(multi14[12][i14]), .B(multi14[13][i14]), .Out(sum14[6][i14]));
      FP16_Add stage032(.A(multi14[14][i14]), .B(multi14[15][i14]), .Out(sum14[7][i14]));
      FP16_Add stage033(.A(multi14[16][i14]), .B(multi14[17][i14]), .Out(sum14[8][i14]));
      FP16_Add stage034(.A(multi14[18][i14]), .B(multi14[19][i14]), .Out(sum14[9][i14]));
      FP16_Add stage035(.A(multi14[20][i14]), .B(multi14[21][i14]), .Out(sum14[10][i14]));
      FP16_Add stage036(.A(multi14[22][i14]), .B(multi14[23][i14]), .Out(sum14[11][i14]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum14[0][i14]), .B(sum14[1][i14]), .Out(sum14[12][i14]));
      FP16_Add stage038(.A(sum14[2][i14]), .B(sum14[3][i14]), .Out(sum14[13][i14]));
      FP16_Add stage039(.A(sum14[4][i14]), .B(sum14[5][i14]), .Out(sum14[14][i14]));
      FP16_Add stage040(.A(sum14[6][i14]), .B(sum14[7][i14]), .Out(sum14[15][i14]));
      FP16_Add stage041(.A(sum14[8][i14]), .B(sum14[9][i14]), .Out(sum14[16][i14]));
      FP16_Add stage042(.A(sum14[10][i14]), .B(sum14[11][i14]), .Out(sum14[17][i14]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum14[12][i14]), .B(sum14[13][i14]), .Out(sum14[18][i14]));
      FP16_Add stage044(.A(sum14[14][i14]), .B(sum14[15][i14]), .Out(sum14[19][i14]));
      FP16_Add stage045(.A(sum14[16][i14]), .B(sum14[17][i14]), .Out(sum14[20][i14]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum14[18][i14]), .B(sum14[19][i14]), .Out(sum14[21][i14]));
      FP16_Add stage047(.A(sum14[20][i14]), .B(multi14[24][i14]), .Out(sum14[22][i14]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum14[21][i14]), .B(sum14[22][i14]), .Out(sum14[23][i14]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum14[23][i14]), .B(feature2Bias), .Out(data_11_array[j14][i14]));
    end
  endgenerate

  ////ROW 15
  generate
    localparam integer j15 = 15;
    for (i15 = 0; i15 < 24; i15 = i15 + 1)
    begin: addbit15
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j15+0][i15+0]), .Out(multi15[0][i15]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j15+0][i15+1]), .Out(multi15[1][i15]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j15+0][i15+2]), .Out(multi15[2][i15]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j15+0][i15+3]), .Out(multi15[3][i15]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j15+0][i15+4]), .Out(multi15[4][i15]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j15+1][i15+0]), .Out(multi15[5][i15]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j15+1][i15+1]), .Out(multi15[6][i15]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j15+1][i15+2]), .Out(multi15[7][i15]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j15+1][i15+3]), .Out(multi15[8][i15]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j15+1][i15+4]), .Out(multi15[9][i15]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j15+2][i15+0]), .Out(multi15[10][i15]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j15+2][i15+1]), .Out(multi15[11][i15]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j15+2][i15+2]), .Out(multi15[12][i15]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j15+2][i15+3]), .Out(multi15[13][i15]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j15+2][i15+4]), .Out(multi15[14][i15]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j15+3][i15+0]), .Out(multi15[15][i15]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j15+3][i15+1]), .Out(multi15[16][i15]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j15+3][i15+2]), .Out(multi15[17][i15]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j15+3][i15+3]), .Out(multi15[18][i15]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j15+3][i15+4]), .Out(multi15[19][i15]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j15+4][i15+0]), .Out(multi15[20][i15]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j15+4][i15+1]), .Out(multi15[21][i15]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j15+4][i15+2]), .Out(multi15[22][i15]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j15+4][i15+3]), .Out(multi15[23][i15]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j15+4][i15+4]), .Out(multi15[24][i15]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi15[0][i15]), .B(multi15[1][i15]), .Out(sum15[0][i15]));
      FP16_Add stage026(.A(multi15[2][i15]), .B(multi15[3][i15]), .Out(sum15[1][i15]));
      FP16_Add stage027(.A(multi15[4][i15]), .B(multi15[5][i15]), .Out(sum15[2][i15]));
      FP16_Add stage028(.A(multi15[6][i15]), .B(multi15[7][i15]), .Out(sum15[3][i15]));
      FP16_Add stage029(.A(multi15[8][i15]), .B(multi15[9][i15]), .Out(sum15[4][i15]));
      FP16_Add stage030(.A(multi15[10][i15]), .B(multi15[11][i15]), .Out(sum15[5][i15]));
      FP16_Add stage031(.A(multi15[12][i15]), .B(multi15[13][i15]), .Out(sum15[6][i15]));
      FP16_Add stage032(.A(multi15[14][i15]), .B(multi15[15][i15]), .Out(sum15[7][i15]));
      FP16_Add stage033(.A(multi15[16][i15]), .B(multi15[17][i15]), .Out(sum15[8][i15]));
      FP16_Add stage034(.A(multi15[18][i15]), .B(multi15[19][i15]), .Out(sum15[9][i15]));
      FP16_Add stage035(.A(multi15[20][i15]), .B(multi15[21][i15]), .Out(sum15[10][i15]));
      FP16_Add stage036(.A(multi15[22][i15]), .B(multi15[23][i15]), .Out(sum15[11][i15]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum15[0][i15]), .B(sum15[1][i15]), .Out(sum15[12][i15]));
      FP16_Add stage038(.A(sum15[2][i15]), .B(sum15[3][i15]), .Out(sum15[13][i15]));
      FP16_Add stage039(.A(sum15[4][i15]), .B(sum15[5][i15]), .Out(sum15[14][i15]));
      FP16_Add stage040(.A(sum15[6][i15]), .B(sum15[7][i15]), .Out(sum15[15][i15]));
      FP16_Add stage041(.A(sum15[8][i15]), .B(sum15[9][i15]), .Out(sum15[16][i15]));
      FP16_Add stage042(.A(sum15[10][i15]), .B(sum15[11][i15]), .Out(sum15[17][i15]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum15[12][i15]), .B(sum15[13][i15]), .Out(sum15[18][i15]));
      FP16_Add stage044(.A(sum15[14][i15]), .B(sum15[15][i15]), .Out(sum15[19][i15]));
      FP16_Add stage045(.A(sum15[16][i15]), .B(sum15[17][i15]), .Out(sum15[20][i15]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum15[18][i15]), .B(sum15[19][i15]), .Out(sum15[21][i15]));
      FP16_Add stage047(.A(sum15[20][i15]), .B(multi15[24][i15]), .Out(sum15[22][i15]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum15[21][i15]), .B(sum15[22][i15]), .Out(sum15[23][i15]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum15[23][i15]), .B(feature2Bias), .Out(data_11_array[j15][i15]));
    end
  endgenerate
  
  ////ROW 16
  generate
    localparam integer j16 = 16;
    for (i16 = 0; i16 < 24; i16 = i16 + 1)
    begin: addbit16
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j16+0][i16+0]), .Out(multi16[0][i16]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j16+0][i16+1]), .Out(multi16[1][i16]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j16+0][i16+2]), .Out(multi16[2][i16]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j16+0][i16+3]), .Out(multi16[3][i16]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j16+0][i16+4]), .Out(multi16[4][i16]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j16+1][i16+0]), .Out(multi16[5][i16]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j16+1][i16+1]), .Out(multi16[6][i16]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j16+1][i16+2]), .Out(multi16[7][i16]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j16+1][i16+3]), .Out(multi16[8][i16]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j16+1][i16+4]), .Out(multi16[9][i16]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j16+2][i16+0]), .Out(multi16[10][i16]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j16+2][i16+1]), .Out(multi16[11][i16]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j16+2][i16+2]), .Out(multi16[12][i16]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j16+2][i16+3]), .Out(multi16[13][i16]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j16+2][i16+4]), .Out(multi16[14][i16]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j16+3][i16+0]), .Out(multi16[15][i16]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j16+3][i16+1]), .Out(multi16[16][i16]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j16+3][i16+2]), .Out(multi16[17][i16]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j16+3][i16+3]), .Out(multi16[18][i16]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j16+3][i16+4]), .Out(multi16[19][i16]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j16+4][i16+0]), .Out(multi16[20][i16]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j16+4][i16+1]), .Out(multi16[21][i16]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j16+4][i16+2]), .Out(multi16[22][i16]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j16+4][i16+3]), .Out(multi16[23][i16]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j16+4][i16+4]), .Out(multi16[24][i16]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi16[0][i16]), .B(multi16[1][i16]), .Out(sum16[0][i16]));
      FP16_Add stage026(.A(multi16[2][i16]), .B(multi16[3][i16]), .Out(sum16[1][i16]));
      FP16_Add stage027(.A(multi16[4][i16]), .B(multi16[5][i16]), .Out(sum16[2][i16]));
      FP16_Add stage028(.A(multi16[6][i16]), .B(multi16[7][i16]), .Out(sum16[3][i16]));
      FP16_Add stage029(.A(multi16[8][i16]), .B(multi16[9][i16]), .Out(sum16[4][i16]));
      FP16_Add stage030(.A(multi16[10][i16]), .B(multi16[11][i16]), .Out(sum16[5][i16]));
      FP16_Add stage031(.A(multi16[12][i16]), .B(multi16[13][i16]), .Out(sum16[6][i16]));
      FP16_Add stage032(.A(multi16[14][i16]), .B(multi16[15][i16]), .Out(sum16[7][i16]));
      FP16_Add stage033(.A(multi16[16][i16]), .B(multi16[17][i16]), .Out(sum16[8][i16]));
      FP16_Add stage034(.A(multi16[18][i16]), .B(multi16[19][i16]), .Out(sum16[9][i16]));
      FP16_Add stage035(.A(multi16[20][i16]), .B(multi16[21][i16]), .Out(sum16[10][i16]));
      FP16_Add stage036(.A(multi16[22][i16]), .B(multi16[23][i16]), .Out(sum16[11][i16]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum16[0][i16]), .B(sum16[1][i16]), .Out(sum16[12][i16]));
      FP16_Add stage038(.A(sum16[2][i16]), .B(sum16[3][i16]), .Out(sum16[13][i16]));
      FP16_Add stage039(.A(sum16[4][i16]), .B(sum16[5][i16]), .Out(sum16[14][i16]));
      FP16_Add stage040(.A(sum16[6][i16]), .B(sum16[7][i16]), .Out(sum16[15][i16]));
      FP16_Add stage041(.A(sum16[8][i16]), .B(sum16[9][i16]), .Out(sum16[16][i16]));
      FP16_Add stage042(.A(sum16[10][i16]), .B(sum16[11][i16]), .Out(sum16[17][i16]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum16[12][i16]), .B(sum16[13][i16]), .Out(sum16[18][i16]));
      FP16_Add stage044(.A(sum16[14][i16]), .B(sum16[15][i16]), .Out(sum16[19][i16]));
      FP16_Add stage045(.A(sum16[16][i16]), .B(sum16[17][i16]), .Out(sum16[20][i16]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum16[18][i16]), .B(sum16[19][i16]), .Out(sum16[21][i16]));
      FP16_Add stage047(.A(sum16[20][i16]), .B(multi16[24][i16]), .Out(sum16[22][i16]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum16[21][i16]), .B(sum16[22][i16]), .Out(sum16[23][i16]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum16[23][i16]), .B(feature2Bias), .Out(data_11_array[j16][i16]));
    end
  endgenerate
  
  ////ROW 17
  generate
    localparam integer j17 = 17;
    for (i17 = 0; i17 < 24; i17 = i17 + 1)
    begin: addbit17
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j17+0][i17+0]), .Out(multi17[0][i17]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j17+0][i17+1]), .Out(multi17[1][i17]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j17+0][i17+2]), .Out(multi17[2][i17]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j17+0][i17+3]), .Out(multi17[3][i17]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j17+0][i17+4]), .Out(multi17[4][i17]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j17+1][i17+0]), .Out(multi17[5][i17]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j17+1][i17+1]), .Out(multi17[6][i17]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j17+1][i17+2]), .Out(multi17[7][i17]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j17+1][i17+3]), .Out(multi17[8][i17]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j17+1][i17+4]), .Out(multi17[9][i17]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j17+2][i17+0]), .Out(multi17[10][i17]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j17+2][i17+1]), .Out(multi17[11][i17]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j17+2][i17+2]), .Out(multi17[12][i17]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j17+2][i17+3]), .Out(multi17[13][i17]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j17+2][i17+4]), .Out(multi17[14][i17]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j17+3][i17+0]), .Out(multi17[15][i17]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j17+3][i17+1]), .Out(multi17[16][i17]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j17+3][i17+2]), .Out(multi17[17][i17]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j17+3][i17+3]), .Out(multi17[18][i17]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j17+3][i17+4]), .Out(multi17[19][i17]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j17+4][i17+0]), .Out(multi17[20][i17]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j17+4][i17+1]), .Out(multi17[21][i17]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j17+4][i17+2]), .Out(multi17[22][i17]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j17+4][i17+3]), .Out(multi17[23][i17]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j17+4][i17+4]), .Out(multi17[24][i17]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi17[0][i17]), .B(multi17[1][i17]), .Out(sum17[0][i17]));
      FP16_Add stage026(.A(multi17[2][i17]), .B(multi17[3][i17]), .Out(sum17[1][i17]));
      FP16_Add stage027(.A(multi17[4][i17]), .B(multi17[5][i17]), .Out(sum17[2][i17]));
      FP16_Add stage028(.A(multi17[6][i17]), .B(multi17[7][i17]), .Out(sum17[3][i17]));
      FP16_Add stage029(.A(multi17[8][i17]), .B(multi17[9][i17]), .Out(sum17[4][i17]));
      FP16_Add stage030(.A(multi17[10][i17]), .B(multi17[11][i17]), .Out(sum17[5][i17]));
      FP16_Add stage031(.A(multi17[12][i17]), .B(multi17[13][i17]), .Out(sum17[6][i17]));
      FP16_Add stage032(.A(multi17[14][i17]), .B(multi17[15][i17]), .Out(sum17[7][i17]));
      FP16_Add stage033(.A(multi17[16][i17]), .B(multi17[17][i17]), .Out(sum17[8][i17]));
      FP16_Add stage034(.A(multi17[18][i17]), .B(multi17[19][i17]), .Out(sum17[9][i17]));
      FP16_Add stage035(.A(multi17[20][i17]), .B(multi17[21][i17]), .Out(sum17[10][i17]));
      FP16_Add stage036(.A(multi17[22][i17]), .B(multi17[23][i17]), .Out(sum17[11][i17]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum17[0][i17]), .B(sum17[1][i17]), .Out(sum17[12][i17]));
      FP16_Add stage038(.A(sum17[2][i17]), .B(sum17[3][i17]), .Out(sum17[13][i17]));
      FP16_Add stage039(.A(sum17[4][i17]), .B(sum17[5][i17]), .Out(sum17[14][i17]));
      FP16_Add stage040(.A(sum17[6][i17]), .B(sum17[7][i17]), .Out(sum17[15][i17]));
      FP16_Add stage041(.A(sum17[8][i17]), .B(sum17[9][i17]), .Out(sum17[16][i17]));
      FP16_Add stage042(.A(sum17[10][i17]), .B(sum17[11][i17]), .Out(sum17[17][i17]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum17[12][i17]), .B(sum17[13][i17]), .Out(sum17[18][i17]));
      FP16_Add stage044(.A(sum17[14][i17]), .B(sum17[15][i17]), .Out(sum17[19][i17]));
      FP16_Add stage045(.A(sum17[16][i17]), .B(sum17[17][i17]), .Out(sum17[20][i17]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum17[18][i17]), .B(sum17[19][i17]), .Out(sum17[21][i17]));
      FP16_Add stage047(.A(sum17[20][i17]), .B(multi17[24][i17]), .Out(sum17[22][i17]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum17[21][i17]), .B(sum17[22][i17]), .Out(sum17[23][i17]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum17[23][i17]), .B(feature2Bias), .Out(data_11_array[j17][i17]));
    end
  endgenerate

////ROW 18
  generate
    localparam integer j18 = 18;
    for (i18 = 0; i18 < 24; i18 = i18 + 1)
    begin: addbit18
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j18+0][i18+0]), .Out(multi18[0][i18]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j18+0][i18+1]), .Out(multi18[1][i18]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j18+0][i18+2]), .Out(multi18[2][i18]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j18+0][i18+3]), .Out(multi18[3][i18]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j18+0][i18+4]), .Out(multi18[4][i18]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j18+1][i18+0]), .Out(multi18[5][i18]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j18+1][i18+1]), .Out(multi18[6][i18]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j18+1][i18+2]), .Out(multi18[7][i18]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j18+1][i18+3]), .Out(multi18[8][i18]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j18+1][i18+4]), .Out(multi18[9][i18]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j18+2][i18+0]), .Out(multi18[10][i18]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j18+2][i18+1]), .Out(multi18[11][i18]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j18+2][i18+2]), .Out(multi18[12][i18]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j18+2][i18+3]), .Out(multi18[13][i18]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j18+2][i18+4]), .Out(multi18[14][i18]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j18+3][i18+0]), .Out(multi18[15][i18]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j18+3][i18+1]), .Out(multi18[16][i18]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j18+3][i18+2]), .Out(multi18[17][i18]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j18+3][i18+3]), .Out(multi18[18][i18]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j18+3][i18+4]), .Out(multi18[19][i18]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j18+4][i18+0]), .Out(multi18[20][i18]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j18+4][i18+1]), .Out(multi18[21][i18]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j18+4][i18+2]), .Out(multi18[22][i18]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j18+4][i18+3]), .Out(multi18[23][i18]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j18+4][i18+4]), .Out(multi18[24][i18]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi18[0][i18]), .B(multi18[1][i18]), .Out(sum18[0][i18]));
      FP16_Add stage026(.A(multi18[2][i18]), .B(multi18[3][i18]), .Out(sum18[1][i18]));
      FP16_Add stage027(.A(multi18[4][i18]), .B(multi18[5][i18]), .Out(sum18[2][i18]));
      FP16_Add stage028(.A(multi18[6][i18]), .B(multi18[7][i18]), .Out(sum18[3][i18]));
      FP16_Add stage029(.A(multi18[8][i18]), .B(multi18[9][i18]), .Out(sum18[4][i18]));
      FP16_Add stage030(.A(multi18[10][i18]), .B(multi18[11][i18]), .Out(sum18[5][i18]));
      FP16_Add stage031(.A(multi18[12][i18]), .B(multi18[13][i18]), .Out(sum18[6][i18]));
      FP16_Add stage032(.A(multi18[14][i18]), .B(multi18[15][i18]), .Out(sum18[7][i18]));
      FP16_Add stage033(.A(multi18[16][i18]), .B(multi18[17][i18]), .Out(sum18[8][i18]));
      FP16_Add stage034(.A(multi18[18][i18]), .B(multi18[19][i18]), .Out(sum18[9][i18]));
      FP16_Add stage035(.A(multi18[20][i18]), .B(multi18[21][i18]), .Out(sum18[10][i18]));
      FP16_Add stage036(.A(multi18[22][i18]), .B(multi18[23][i18]), .Out(sum18[11][i18]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum18[0][i18]), .B(sum18[1][i18]), .Out(sum18[12][i18]));
      FP16_Add stage038(.A(sum18[2][i18]), .B(sum18[3][i18]), .Out(sum18[13][i18]));
      FP16_Add stage039(.A(sum18[4][i18]), .B(sum18[5][i18]), .Out(sum18[14][i18]));
      FP16_Add stage040(.A(sum18[6][i18]), .B(sum18[7][i18]), .Out(sum18[15][i18]));
      FP16_Add stage041(.A(sum18[8][i18]), .B(sum18[9][i18]), .Out(sum18[16][i18]));
      FP16_Add stage042(.A(sum18[10][i18]), .B(sum18[11][i18]), .Out(sum18[17][i18]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum18[12][i18]), .B(sum18[13][i18]), .Out(sum18[18][i18]));
      FP16_Add stage044(.A(sum18[14][i18]), .B(sum18[15][i18]), .Out(sum18[19][i18]));
      FP16_Add stage045(.A(sum18[16][i18]), .B(sum18[17][i18]), .Out(sum18[20][i18]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum18[18][i18]), .B(sum18[19][i18]), .Out(sum18[21][i18]));
      FP16_Add stage047(.A(sum18[20][i18]), .B(multi18[24][i18]), .Out(sum18[22][i18]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum18[21][i18]), .B(sum18[22][i18]), .Out(sum18[23][i18]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum18[23][i18]), .B(feature2Bias), .Out(data_11_array[j18][i18]));
    end
  endgenerate

////ROW 19
  generate
    localparam integer j19 = 19;
    for (i19 = 0; i19 < 24; i19 = i19 + 1)
    begin: addbit19
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j19+0][i19+0]), .Out(multi19[0][i19]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j19+0][i19+1]), .Out(multi19[1][i19]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j19+0][i19+2]), .Out(multi19[2][i19]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j19+0][i19+3]), .Out(multi19[3][i19]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j19+0][i19+4]), .Out(multi19[4][i19]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j19+1][i19+0]), .Out(multi19[5][i19]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j19+1][i19+1]), .Out(multi19[6][i19]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j19+1][i19+2]), .Out(multi19[7][i19]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j19+1][i19+3]), .Out(multi19[8][i19]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j19+1][i19+4]), .Out(multi19[9][i19]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j19+2][i19+0]), .Out(multi19[10][i19]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j19+2][i19+1]), .Out(multi19[11][i19]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j19+2][i19+2]), .Out(multi19[12][i19]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j19+2][i19+3]), .Out(multi19[13][i19]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j19+2][i19+4]), .Out(multi19[14][i19]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j19+3][i19+0]), .Out(multi19[15][i19]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j19+3][i19+1]), .Out(multi19[16][i19]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j19+3][i19+2]), .Out(multi19[17][i19]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j19+3][i19+3]), .Out(multi19[18][i19]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j19+3][i19+4]), .Out(multi19[19][i19]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j19+4][i19+0]), .Out(multi19[20][i19]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j19+4][i19+1]), .Out(multi19[21][i19]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j19+4][i19+2]), .Out(multi19[22][i19]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j19+4][i19+3]), .Out(multi19[23][i19]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j19+4][i19+4]), .Out(multi19[24][i19]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi19[0][i19]), .B(multi19[1][i19]), .Out(sum19[0][i19]));
      FP16_Add stage026(.A(multi19[2][i19]), .B(multi19[3][i19]), .Out(sum19[1][i19]));
      FP16_Add stage027(.A(multi19[4][i19]), .B(multi19[5][i19]), .Out(sum19[2][i19]));
      FP16_Add stage028(.A(multi19[6][i19]), .B(multi19[7][i19]), .Out(sum19[3][i19]));
      FP16_Add stage029(.A(multi19[8][i19]), .B(multi19[9][i19]), .Out(sum19[4][i19]));
      FP16_Add stage030(.A(multi19[10][i19]), .B(multi19[11][i19]), .Out(sum19[5][i19]));
      FP16_Add stage031(.A(multi19[12][i19]), .B(multi19[13][i19]), .Out(sum19[6][i19]));
      FP16_Add stage032(.A(multi19[14][i19]), .B(multi19[15][i19]), .Out(sum19[7][i19]));
      FP16_Add stage033(.A(multi19[16][i19]), .B(multi19[17][i19]), .Out(sum19[8][i19]));
      FP16_Add stage034(.A(multi19[18][i19]), .B(multi19[19][i19]), .Out(sum19[9][i19]));
      FP16_Add stage035(.A(multi19[20][i19]), .B(multi19[21][i19]), .Out(sum19[10][i19]));
      FP16_Add stage036(.A(multi19[22][i19]), .B(multi19[23][i19]), .Out(sum19[11][i19]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum19[0][i19]), .B(sum19[1][i19]), .Out(sum19[12][i19]));
      FP16_Add stage038(.A(sum19[2][i19]), .B(sum19[3][i19]), .Out(sum19[13][i19]));
      FP16_Add stage039(.A(sum19[4][i19]), .B(sum19[5][i19]), .Out(sum19[14][i19]));
      FP16_Add stage040(.A(sum19[6][i19]), .B(sum19[7][i19]), .Out(sum19[15][i19]));
      FP16_Add stage041(.A(sum19[8][i19]), .B(sum19[9][i19]), .Out(sum19[16][i19]));
      FP16_Add stage042(.A(sum19[10][i19]), .B(sum19[11][i19]), .Out(sum19[17][i19]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum19[12][i19]), .B(sum19[13][i19]), .Out(sum19[18][i19]));
      FP16_Add stage044(.A(sum19[14][i19]), .B(sum19[15][i19]), .Out(sum19[19][i19]));
      FP16_Add stage045(.A(sum19[16][i19]), .B(sum19[17][i19]), .Out(sum19[20][i19]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum19[18][i19]), .B(sum19[19][i19]), .Out(sum19[21][i19]));
      FP16_Add stage047(.A(sum19[20][i19]), .B(multi19[24][i19]), .Out(sum19[22][i19]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum19[21][i19]), .B(sum19[22][i19]), .Out(sum19[23][i19]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum19[23][i19]), .B(feature2Bias), .Out(data_11_array[j19][i19]));
    end
  endgenerate

////ROW 20
  generate
    localparam integer j20 = 20;
    for (i20 = 0; i20 < 24; i20 = i20 + 1)
    begin: addbit20
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j20+0][i20+0]), .Out(multi20[0][i20]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j20+0][i20+1]), .Out(multi20[1][i20]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j20+0][i20+2]), .Out(multi20[2][i20]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j20+0][i20+3]), .Out(multi20[3][i20]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j20+0][i20+4]), .Out(multi20[4][i20]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j20+1][i20+0]), .Out(multi20[5][i20]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j20+1][i20+1]), .Out(multi20[6][i20]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j20+1][i20+2]), .Out(multi20[7][i20]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j20+1][i20+3]), .Out(multi20[8][i20]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j20+1][i20+4]), .Out(multi20[9][i20]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j20+2][i20+0]), .Out(multi20[10][i20]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j20+2][i20+1]), .Out(multi20[11][i20]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j20+2][i20+2]), .Out(multi20[12][i20]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j20+2][i20+3]), .Out(multi20[13][i20]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j20+2][i20+4]), .Out(multi20[14][i20]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j20+3][i20+0]), .Out(multi20[15][i20]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j20+3][i20+1]), .Out(multi20[16][i20]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j20+3][i20+2]), .Out(multi20[17][i20]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j20+3][i20+3]), .Out(multi20[18][i20]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j20+3][i20+4]), .Out(multi20[19][i20]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j20+4][i20+0]), .Out(multi20[20][i20]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j20+4][i20+1]), .Out(multi20[21][i20]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j20+4][i20+2]), .Out(multi20[22][i20]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j20+4][i20+3]), .Out(multi20[23][i20]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j20+4][i20+4]), .Out(multi20[24][i20]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi20[0][i20]), .B(multi20[1][i20]), .Out(sum20[0][i20]));
      FP16_Add stage026(.A(multi20[2][i20]), .B(multi20[3][i20]), .Out(sum20[1][i20]));
      FP16_Add stage027(.A(multi20[4][i20]), .B(multi20[5][i20]), .Out(sum20[2][i20]));
      FP16_Add stage028(.A(multi20[6][i20]), .B(multi20[7][i20]), .Out(sum20[3][i20]));
      FP16_Add stage029(.A(multi20[8][i20]), .B(multi20[9][i20]), .Out(sum20[4][i20]));
      FP16_Add stage030(.A(multi20[10][i20]), .B(multi20[11][i20]), .Out(sum20[5][i20]));
      FP16_Add stage031(.A(multi20[12][i20]), .B(multi20[13][i20]), .Out(sum20[6][i20]));
      FP16_Add stage032(.A(multi20[14][i20]), .B(multi20[15][i20]), .Out(sum20[7][i20]));
      FP16_Add stage033(.A(multi20[16][i20]), .B(multi20[17][i20]), .Out(sum20[8][i20]));
      FP16_Add stage034(.A(multi20[18][i20]), .B(multi20[19][i20]), .Out(sum20[9][i20]));
      FP16_Add stage035(.A(multi20[20][i20]), .B(multi20[21][i20]), .Out(sum20[10][i20]));
      FP16_Add stage036(.A(multi20[22][i20]), .B(multi20[23][i20]), .Out(sum20[11][i20]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum20[0][i20]), .B(sum20[1][i20]), .Out(sum20[12][i20]));
      FP16_Add stage038(.A(sum20[2][i20]), .B(sum20[3][i20]), .Out(sum20[13][i20]));
      FP16_Add stage039(.A(sum20[4][i20]), .B(sum20[5][i20]), .Out(sum20[14][i20]));
      FP16_Add stage040(.A(sum20[6][i20]), .B(sum20[7][i20]), .Out(sum20[15][i20]));
      FP16_Add stage041(.A(sum20[8][i20]), .B(sum20[9][i20]), .Out(sum20[16][i20]));
      FP16_Add stage042(.A(sum20[10][i20]), .B(sum20[11][i20]), .Out(sum20[17][i20]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum20[12][i20]), .B(sum20[13][i20]), .Out(sum20[18][i20]));
      FP16_Add stage044(.A(sum20[14][i20]), .B(sum20[15][i20]), .Out(sum20[19][i20]));
      FP16_Add stage045(.A(sum20[16][i20]), .B(sum20[17][i20]), .Out(sum20[20][i20]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum20[18][i20]), .B(sum20[19][i20]), .Out(sum20[21][i20]));
      FP16_Add stage047(.A(sum20[20][i20]), .B(multi20[24][i20]), .Out(sum20[22][i20]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum20[21][i20]), .B(sum20[22][i20]), .Out(sum20[23][i20]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum20[23][i20]), .B(feature2Bias), .Out(data_11_array[j20][i20]));
    end
  endgenerate

////ROW 21
  generate
    localparam integer j21 = 21;
    for (i21 = 0; i21 < 24; i21 = i21 + 1)
    begin: addbit21
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j21+0][i21+0]), .Out(multi21[0][i21]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j21+0][i21+1]), .Out(multi21[1][i21]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j21+0][i21+2]), .Out(multi21[2][i21]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j21+0][i21+3]), .Out(multi21[3][i21]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j21+0][i21+4]), .Out(multi21[4][i21]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j21+1][i21+0]), .Out(multi21[5][i21]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j21+1][i21+1]), .Out(multi21[6][i21]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j21+1][i21+2]), .Out(multi21[7][i21]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j21+1][i21+3]), .Out(multi21[8][i21]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j21+1][i21+4]), .Out(multi21[9][i21]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j21+2][i21+0]), .Out(multi21[10][i21]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j21+2][i21+1]), .Out(multi21[11][i21]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j21+2][i21+2]), .Out(multi21[12][i21]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j21+2][i21+3]), .Out(multi21[13][i21]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j21+2][i21+4]), .Out(multi21[14][i21]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j21+3][i21+0]), .Out(multi21[15][i21]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j21+3][i21+1]), .Out(multi21[16][i21]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j21+3][i21+2]), .Out(multi21[17][i21]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j21+3][i21+3]), .Out(multi21[18][i21]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j21+3][i21+4]), .Out(multi21[19][i21]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j21+4][i21+0]), .Out(multi21[20][i21]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j21+4][i21+1]), .Out(multi21[21][i21]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j21+4][i21+2]), .Out(multi21[22][i21]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j21+4][i21+3]), .Out(multi21[23][i21]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j21+4][i21+4]), .Out(multi21[24][i21]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi21[0][i21]), .B(multi21[1][i21]), .Out(sum21[0][i21]));
      FP16_Add stage026(.A(multi21[2][i21]), .B(multi21[3][i21]), .Out(sum21[1][i21]));
      FP16_Add stage027(.A(multi21[4][i21]), .B(multi21[5][i21]), .Out(sum21[2][i21]));
      FP16_Add stage028(.A(multi21[6][i21]), .B(multi21[7][i21]), .Out(sum21[3][i21]));
      FP16_Add stage029(.A(multi21[8][i21]), .B(multi21[9][i21]), .Out(sum21[4][i21]));
      FP16_Add stage030(.A(multi21[10][i21]), .B(multi21[11][i21]), .Out(sum21[5][i21]));
      FP16_Add stage031(.A(multi21[12][i21]), .B(multi21[13][i21]), .Out(sum21[6][i21]));
      FP16_Add stage032(.A(multi21[14][i21]), .B(multi21[15][i21]), .Out(sum21[7][i21]));
      FP16_Add stage033(.A(multi21[16][i21]), .B(multi21[17][i21]), .Out(sum21[8][i21]));
      FP16_Add stage034(.A(multi21[18][i21]), .B(multi21[19][i21]), .Out(sum21[9][i21]));
      FP16_Add stage035(.A(multi21[20][i21]), .B(multi21[21][i21]), .Out(sum21[10][i21]));
      FP16_Add stage036(.A(multi21[22][i21]), .B(multi21[23][i21]), .Out(sum21[11][i21]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum21[0][i21]), .B(sum21[1][i21]), .Out(sum21[12][i21]));
      FP16_Add stage038(.A(sum21[2][i21]), .B(sum21[3][i21]), .Out(sum21[13][i21]));
      FP16_Add stage039(.A(sum21[4][i21]), .B(sum21[5][i21]), .Out(sum21[14][i21]));
      FP16_Add stage040(.A(sum21[6][i21]), .B(sum21[7][i21]), .Out(sum21[15][i21]));
      FP16_Add stage041(.A(sum21[8][i21]), .B(sum21[9][i21]), .Out(sum21[16][i21]));
      FP16_Add stage042(.A(sum21[10][i21]), .B(sum21[11][i21]), .Out(sum21[17][i21]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum21[12][i21]), .B(sum21[13][i21]), .Out(sum21[18][i21]));
      FP16_Add stage044(.A(sum21[14][i21]), .B(sum21[15][i21]), .Out(sum21[19][i21]));
      FP16_Add stage045(.A(sum21[16][i21]), .B(sum21[17][i21]), .Out(sum21[20][i21]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum21[18][i21]), .B(sum21[19][i21]), .Out(sum21[21][i21]));
      FP16_Add stage047(.A(sum21[20][i21]), .B(multi21[24][i21]), .Out(sum21[22][i21]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum21[21][i21]), .B(sum21[22][i21]), .Out(sum21[23][i21]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum21[23][i21]), .B(feature2Bias), .Out(data_11_array[j21][i21]));
    end
  endgenerate

////ROW 22
  generate
    localparam integer j22 = 22;
    for (i22 = 0; i22 < 24; i22 = i22 + 1)
    begin: addbit22
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j22+0][i22+0]), .Out(multi22[0][i22]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j22+0][i22+1]), .Out(multi22[1][i22]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j22+0][i22+2]), .Out(multi22[2][i22]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j22+0][i22+3]), .Out(multi22[3][i22]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j22+0][i22+4]), .Out(multi22[4][i22]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j22+1][i22+0]), .Out(multi22[5][i22]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j22+1][i22+1]), .Out(multi22[6][i22]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j22+1][i22+2]), .Out(multi22[7][i22]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j22+1][i22+3]), .Out(multi22[8][i22]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j22+1][i22+4]), .Out(multi22[9][i22]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j22+2][i22+0]), .Out(multi22[10][i22]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j22+2][i22+1]), .Out(multi22[11][i22]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j22+2][i22+2]), .Out(multi22[12][i22]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j22+2][i22+3]), .Out(multi22[13][i22]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j22+2][i22+4]), .Out(multi22[14][i22]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j22+3][i22+0]), .Out(multi22[15][i22]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j22+3][i22+1]), .Out(multi22[16][i22]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j22+3][i22+2]), .Out(multi22[17][i22]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j22+3][i22+3]), .Out(multi22[18][i22]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j22+3][i22+4]), .Out(multi22[19][i22]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j22+4][i22+0]), .Out(multi22[20][i22]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j22+4][i22+1]), .Out(multi22[21][i22]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j22+4][i22+2]), .Out(multi22[22][i22]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j22+4][i22+3]), .Out(multi22[23][i22]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j22+4][i22+4]), .Out(multi22[24][i22]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi22[0][i22]), .B(multi22[1][i22]), .Out(sum22[0][i22]));
      FP16_Add stage026(.A(multi22[2][i22]), .B(multi22[3][i22]), .Out(sum22[1][i22]));
      FP16_Add stage027(.A(multi22[4][i22]), .B(multi22[5][i22]), .Out(sum22[2][i22]));
      FP16_Add stage028(.A(multi22[6][i22]), .B(multi22[7][i22]), .Out(sum22[3][i22]));
      FP16_Add stage029(.A(multi22[8][i22]), .B(multi22[9][i22]), .Out(sum22[4][i22]));
      FP16_Add stage030(.A(multi22[10][i22]), .B(multi22[11][i22]), .Out(sum22[5][i22]));
      FP16_Add stage031(.A(multi22[12][i22]), .B(multi22[13][i22]), .Out(sum22[6][i22]));
      FP16_Add stage032(.A(multi22[14][i22]), .B(multi22[15][i22]), .Out(sum22[7][i22]));
      FP16_Add stage033(.A(multi22[16][i22]), .B(multi22[17][i22]), .Out(sum22[8][i22]));
      FP16_Add stage034(.A(multi22[18][i22]), .B(multi22[19][i22]), .Out(sum22[9][i22]));
      FP16_Add stage035(.A(multi22[20][i22]), .B(multi22[21][i22]), .Out(sum22[10][i22]));
      FP16_Add stage036(.A(multi22[22][i22]), .B(multi22[23][i22]), .Out(sum22[11][i22]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum22[0][i22]), .B(sum22[1][i22]), .Out(sum22[12][i22]));
      FP16_Add stage038(.A(sum22[2][i22]), .B(sum22[3][i22]), .Out(sum22[13][i22]));
      FP16_Add stage039(.A(sum22[4][i22]), .B(sum22[5][i22]), .Out(sum22[14][i22]));
      FP16_Add stage040(.A(sum22[6][i22]), .B(sum22[7][i22]), .Out(sum22[15][i22]));
      FP16_Add stage041(.A(sum22[8][i22]), .B(sum22[9][i22]), .Out(sum22[16][i22]));
      FP16_Add stage042(.A(sum22[10][i22]), .B(sum22[11][i22]), .Out(sum22[17][i22]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum22[12][i22]), .B(sum22[13][i22]), .Out(sum22[18][i22]));
      FP16_Add stage044(.A(sum22[14][i22]), .B(sum22[15][i22]), .Out(sum22[19][i22]));
      FP16_Add stage045(.A(sum22[16][i22]), .B(sum22[17][i22]), .Out(sum22[20][i22]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum22[18][i22]), .B(sum22[19][i22]), .Out(sum22[21][i22]));
      FP16_Add stage047(.A(sum22[20][i22]), .B(multi22[24][i22]), .Out(sum22[22][i22]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum22[21][i22]), .B(sum22[22][i22]), .Out(sum22[23][i22]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum22[23][i22]), .B(feature2Bias), .Out(data_11_array[j22][i22]));
    end
  endgenerate

////ROW 23
  generate
    localparam integer j23 = 23;
    for (i23 = 0; i23 < 24; i23 = i23 + 1)
    begin: addbit23
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j23+0][i23+0]), .Out(multi23[0][i23]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j23+0][i23+1]), .Out(multi23[1][i23]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j23+0][i23+2]), .Out(multi23[2][i23]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j23+0][i23+3]), .Out(multi23[3][i23]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j23+0][i23+4]), .Out(multi23[4][i23]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j23+1][i23+0]), .Out(multi23[5][i23]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j23+1][i23+1]), .Out(multi23[6][i23]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j23+1][i23+2]), .Out(multi23[7][i23]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j23+1][i23+3]), .Out(multi23[8][i23]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j23+1][i23+4]), .Out(multi23[9][i23]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j23+2][i23+0]), .Out(multi23[10][i23]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j23+2][i23+1]), .Out(multi23[11][i23]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j23+2][i23+2]), .Out(multi23[12][i23]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j23+2][i23+3]), .Out(multi23[13][i23]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j23+2][i23+4]), .Out(multi23[14][i23]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j23+3][i23+0]), .Out(multi23[15][i23]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j23+3][i23+1]), .Out(multi23[16][i23]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j23+3][i23+2]), .Out(multi23[17][i23]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j23+3][i23+3]), .Out(multi23[18][i23]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j23+3][i23+4]), .Out(multi23[19][i23]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j23+4][i23+0]), .Out(multi23[20][i23]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j23+4][i23+1]), .Out(multi23[21][i23]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j23+4][i23+2]), .Out(multi23[22][i23]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j23+4][i23+3]), .Out(multi23[23][i23]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j23+4][i23+4]), .Out(multi23[24][i23]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi23[0][i23]), .B(multi23[1][i23]), .Out(sum23[0][i23]));
      FP16_Add stage026(.A(multi23[2][i23]), .B(multi23[3][i23]), .Out(sum23[1][i23]));
      FP16_Add stage027(.A(multi23[4][i23]), .B(multi23[5][i23]), .Out(sum23[2][i23]));
      FP16_Add stage028(.A(multi23[6][i23]), .B(multi23[7][i23]), .Out(sum23[3][i23]));
      FP16_Add stage029(.A(multi23[8][i23]), .B(multi23[9][i23]), .Out(sum23[4][i23]));
      FP16_Add stage030(.A(multi23[10][i23]), .B(multi23[11][i23]), .Out(sum23[5][i23]));
      FP16_Add stage031(.A(multi23[12][i23]), .B(multi23[13][i23]), .Out(sum23[6][i23]));
      FP16_Add stage032(.A(multi23[14][i23]), .B(multi23[15][i23]), .Out(sum23[7][i23]));
      FP16_Add stage033(.A(multi23[16][i23]), .B(multi23[17][i23]), .Out(sum23[8][i23]));
      FP16_Add stage034(.A(multi23[18][i23]), .B(multi23[19][i23]), .Out(sum23[9][i23]));
      FP16_Add stage035(.A(multi23[20][i23]), .B(multi23[21][i23]), .Out(sum23[10][i23]));
      FP16_Add stage036(.A(multi23[22][i23]), .B(multi23[23][i23]), .Out(sum23[11][i23]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum23[0][i23]), .B(sum23[1][i23]), .Out(sum23[12][i23]));
      FP16_Add stage038(.A(sum23[2][i23]), .B(sum23[3][i23]), .Out(sum23[13][i23]));
      FP16_Add stage039(.A(sum23[4][i23]), .B(sum23[5][i23]), .Out(sum23[14][i23]));
      FP16_Add stage040(.A(sum23[6][i23]), .B(sum23[7][i23]), .Out(sum23[15][i23]));
      FP16_Add stage041(.A(sum23[8][i23]), .B(sum23[9][i23]), .Out(sum23[16][i23]));
      FP16_Add stage042(.A(sum23[10][i23]), .B(sum23[11][i23]), .Out(sum23[17][i23]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum23[12][i23]), .B(sum23[13][i23]), .Out(sum23[18][i23]));
      FP16_Add stage044(.A(sum23[14][i23]), .B(sum23[15][i23]), .Out(sum23[19][i23]));
      FP16_Add stage045(.A(sum23[16][i23]), .B(sum23[17][i23]), .Out(sum23[20][i23]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum23[18][i23]), .B(sum23[19][i23]), .Out(sum23[21][i23]));
      FP16_Add stage047(.A(sum23[20][i23]), .B(multi23[24][i23]), .Out(sum23[22][i23]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum23[21][i23]), .B(sum23[22][i23]), .Out(sum23[23][i23]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum23[23][i23]), .B(feature2Bias), .Out(data_11_array[j23][i23]));
    end
  endgenerate

////ROW 24
  generate
    localparam integer j24 = 24;
    for (i24 = 0; i24 < 24; i24 = i24 + 1)
    begin: addbit24
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature2Weight_0), .B(data_array[j24+0][i24+0]), .Out(multi24[0][i24]));
      FP16_Multiply stage01(.A(feature2Weight_1), .B(data_array[j24+0][i24+1]), .Out(multi24[1][i24]));
      FP16_Multiply stage02(.A(feature2Weight_2), .B(data_array[j24+0][i24+2]), .Out(multi24[2][i24]));
      FP16_Multiply stage03(.A(feature2Weight_3), .B(data_array[j24+0][i24+3]), .Out(multi24[3][i24]));
      FP16_Multiply stage04(.A(feature2Weight_4), .B(data_array[j24+0][i24+4]), .Out(multi24[4][i24]));
      FP16_Multiply stage05(.A(feature2Weight_5), .B(data_array[j24+1][i24+0]), .Out(multi24[5][i24]));
      FP16_Multiply stage06(.A(feature2Weight_6), .B(data_array[j24+1][i24+1]), .Out(multi24[6][i24]));
      FP16_Multiply stage07(.A(feature2Weight_7), .B(data_array[j24+1][i24+2]), .Out(multi24[7][i24]));
      FP16_Multiply stage08(.A(feature2Weight_8), .B(data_array[j24+1][i24+3]), .Out(multi24[8][i24]));
      FP16_Multiply stage09(.A(feature2Weight_9), .B(data_array[j24+1][i24+4]), .Out(multi24[9][i24]));
      FP16_Multiply stage010(.A(feature2Weight_10), .B(data_array[j24+2][i24+0]), .Out(multi24[10][i24]));
      FP16_Multiply stage011(.A(feature2Weight_11), .B(data_array[j24+2][i24+1]), .Out(multi24[11][i24]));
      FP16_Multiply stage012(.A(feature2Weight_12), .B(data_array[j24+2][i24+2]), .Out(multi24[12][i24]));
      FP16_Multiply stage013(.A(feature2Weight_13), .B(data_array[j24+2][i24+3]), .Out(multi24[13][i24]));
      FP16_Multiply stage014(.A(feature2Weight_14), .B(data_array[j24+2][i24+4]), .Out(multi24[14][i24]));
      FP16_Multiply stage015(.A(feature2Weight_15), .B(data_array[j24+3][i24+0]), .Out(multi24[15][i24]));
      FP16_Multiply stage016(.A(feature2Weight_16), .B(data_array[j24+3][i24+1]), .Out(multi24[16][i24]));
      FP16_Multiply stage017(.A(feature2Weight_17), .B(data_array[j24+3][i24+2]), .Out(multi24[17][i24]));
      FP16_Multiply stage018(.A(feature2Weight_18), .B(data_array[j24+3][i24+3]), .Out(multi24[18][i24]));
      FP16_Multiply stage019(.A(feature2Weight_19), .B(data_array[j24+3][i24+4]), .Out(multi24[19][i24]));
      FP16_Multiply stage020(.A(feature2Weight_20), .B(data_array[j24+4][i24+0]), .Out(multi24[20][i24]));
      FP16_Multiply stage021(.A(feature2Weight_21), .B(data_array[j24+4][i24+1]), .Out(multi24[21][i24]));
      FP16_Multiply stage022(.A(feature2Weight_22), .B(data_array[j24+4][i24+2]), .Out(multi24[22][i24]));
      FP16_Multiply stage023(.A(feature2Weight_23), .B(data_array[j24+4][i24+3]), .Out(multi24[23][i24]));
      FP16_Multiply stage024(.A(feature2Weight_24), .B(data_array[j24+4][i24+4]), .Out(multi24[24][i24]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi24[0][i24]), .B(multi24[1][i24]), .Out(sum24[0][i24]));
      FP16_Add stage026(.A(multi24[2][i24]), .B(multi24[3][i24]), .Out(sum24[1][i24]));
      FP16_Add stage027(.A(multi24[4][i24]), .B(multi24[5][i24]), .Out(sum24[2][i24]));
      FP16_Add stage028(.A(multi24[6][i24]), .B(multi24[7][i24]), .Out(sum24[3][i24]));
      FP16_Add stage029(.A(multi24[8][i24]), .B(multi24[9][i24]), .Out(sum24[4][i24]));
      FP16_Add stage030(.A(multi24[10][i24]), .B(multi24[11][i24]), .Out(sum24[5][i24]));
      FP16_Add stage031(.A(multi24[12][i24]), .B(multi24[13][i24]), .Out(sum24[6][i24]));
      FP16_Add stage032(.A(multi24[14][i24]), .B(multi24[15][i24]), .Out(sum24[7][i24]));
      FP16_Add stage033(.A(multi24[16][i24]), .B(multi24[17][i24]), .Out(sum24[8][i24]));
      FP16_Add stage034(.A(multi24[18][i24]), .B(multi24[19][i24]), .Out(sum24[9][i24]));
      FP16_Add stage035(.A(multi24[20][i24]), .B(multi24[21][i24]), .Out(sum24[10][i24]));
      FP16_Add stage036(.A(multi24[22][i24]), .B(multi24[23][i24]), .Out(sum24[11][i24]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum24[0][i24]), .B(sum24[1][i24]), .Out(sum24[12][i24]));
      FP16_Add stage038(.A(sum24[2][i24]), .B(sum24[3][i24]), .Out(sum24[13][i24]));
      FP16_Add stage039(.A(sum24[4][i24]), .B(sum24[5][i24]), .Out(sum24[14][i24]));
      FP16_Add stage040(.A(sum24[6][i24]), .B(sum24[7][i24]), .Out(sum24[15][i24]));
      FP16_Add stage041(.A(sum24[8][i24]), .B(sum24[9][i24]), .Out(sum24[16][i24]));
      FP16_Add stage042(.A(sum24[10][i24]), .B(sum24[11][i24]), .Out(sum24[17][i24]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum24[12][i24]), .B(sum24[13][i24]), .Out(sum24[18][i24]));
      FP16_Add stage044(.A(sum24[14][i24]), .B(sum24[15][i24]), .Out(sum24[19][i24]));
      FP16_Add stage045(.A(sum24[16][i24]), .B(sum24[17][i24]), .Out(sum24[20][i24]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum24[18][i24]), .B(sum24[19][i24]), .Out(sum24[21][i24]));
      FP16_Add stage047(.A(sum24[20][i24]), .B(multi24[24][i24]), .Out(sum24[22][i24]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum24[21][i24]), .B(sum24[22][i24]), .Out(sum24[23][i24]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum24[23][i24]), .B(feature2Bias), .Out(data_11_array[j24][i24]));
    end
  endgenerate
  
  localparam integer c0 = 0;
    generate 
        localparam integer d0 = 0;
        for (n0 = 0; n0 < 16; n0 = n0 + 1) 
        begin: outbit0
            assign data_11[n0 + d0*16 + c0*28*16] = data_11_array[c0][d0][n0];
        end
    endgenerate
    generate 
        localparam integer d1 = 1;
        for (n1 = 0; n1 < 16; n1 = n1 + 1) 
        begin: outbit1
            assign data_11[n1 + d1*16 + c0*28*16] = data_11_array[c0][d1][n1];
        end
    endgenerate
    generate 
        localparam integer d2 = 2;
        for (n2 = 0; n2 < 16; n2 = n2 + 1) 
        begin: outbit2
            assign data_11[n2 + d2*16 + c0*28*16] = data_11_array[c0][d2][n2];
        end
    endgenerate
    generate 
        localparam integer d3 = 3;
        for (n3 = 0; n3 < 16; n3 = n3 + 1) 
        begin: outbit3
            assign data_11[n3 + d3*16 + c0*28*16] = data_11_array[c0][d3][n3];
        end
    endgenerate
    generate 
        localparam integer d4 = 4;
        for (n4 = 0; n4 < 16; n4 = n4 + 1) 
        begin: outbit4
            assign data_11[n4 + d4*16 + c0*28*16] = data_11_array[c0][d4][n4];
        end
    endgenerate
    generate 
        localparam integer d5 = 5;
        for (n5 = 0; n5 < 16; n5 = n5 + 1) 
        begin: outbit5
            assign data_11[n5 + d5*16 + c0*28*16] = data_11_array[c0][d5][n5];
        end
    endgenerate
    generate 
        localparam integer d6 = 6;
        for (n6 = 0; n6 < 16; n6 = n6 + 1) 
        begin: outbit6
            assign data_11[n6 + d6*16 + c0*28*16] = data_11_array[c0][d6][n6];
        end
    endgenerate
    generate 
        localparam integer d7 = 7;
        for (n7 = 0; n7 < 16; n7 = n7 + 1) 
        begin: outbit7
            assign data_11[n7 + d7*16 + c0*28*16] = data_11_array[c0][d7][n7];
        end
    endgenerate
    generate 
        localparam integer d8 = 8;
        for (n8 = 0; n8 < 16; n8 = n8 + 1) 
        begin: outbit8
            assign data_11[n8 + d8*16 + c0*28*16] = data_11_array[c0][d8][n8];
        end
    endgenerate
    generate 
        localparam integer d9 = 9;
        for (n9 = 0; n9 < 16; n9 = n9 + 1) 
        begin: outbit9
            assign data_11[n9 + d9*16 + c0*28*16] = data_11_array[c0][d9][n9];
        end
    endgenerate
    generate 
        localparam integer d10 = 10;
        for (n10 = 0; n10 < 16; n10 = n10 + 1) 
        begin: outbit10
            assign data_11[n10 + d10*16 + c0*28*16] = data_11_array[c0][d10][n10];
        end
    endgenerate
    generate 
        localparam integer d11 = 11;
        for (n11 = 0; n11 < 16; n11 = n11 + 1) 
        begin: outbit11
            assign data_11[n11 + d11*16 + c0*28*16] = data_11_array[c0][d11][n11];
        end
    endgenerate
    generate 
        localparam integer d12 = 12;
        for (n12 = 0; n12 < 16; n12 = n12 + 1) 
        begin: outbit12
            assign data_11[n12 + d12*16 + c0*28*16] = data_11_array[c0][d12][n12];
        end
    endgenerate
    generate 
        localparam integer d13 = 13;
        for (n13 = 0; n13 < 16; n13 = n13 + 1) 
        begin: outbit13
            assign data_11[n13 + d13*16 + c0*28*16] = data_11_array[c0][d13][n13];
        end
    endgenerate
    generate 
        localparam integer d14 = 14;
        for (n14 = 0; n14 < 16; n14 = n14 + 1) 
        begin: outbit14
            assign data_11[n14 + d14*16 + c0*28*16] = data_11_array[c0][d14][n14];
        end
    endgenerate
    generate 
        localparam integer d15 = 15;
        for (n15 = 0; n15 < 16; n15 = n15 + 1) 
        begin: outbit15
            assign data_11[n15 + d15*16 + c0*28*16] = data_11_array[c0][d15][n15];
        end
    endgenerate
    generate 
        localparam integer d16 = 16;
        for (n16 = 0; n16 < 16; n16 = n16 + 1) 
        begin: outbit16
            assign data_11[n16 + d16*16 + c0*28*16] = data_11_array[c0][d16][n16];
        end
    endgenerate
    generate 
        localparam integer d17 = 17;
        for (n17 = 0; n17 < 16; n17 = n17 + 1) 
        begin: outbit17
            assign data_11[n17 + d17*16 + c0*28*16] = data_11_array[c0][d17][n17];
        end
    endgenerate
    generate 
        localparam integer d18 = 18;
        for (n18 = 0; n18 < 16; n18 = n18 + 1) 
        begin: outbit18
            assign data_11[n18 + d18*16 + c0*28*16] = data_11_array[c0][d18][n18];
        end
    endgenerate
    generate 
        localparam integer d19 = 19;
        for (n19 = 0; n19 < 16; n19 = n19 + 1) 
        begin: outbit19
            assign data_11[n19 + d19*16 + c0*28*16] = data_11_array[c0][d19][n19];
        end
    endgenerate
    generate 
        localparam integer d20 = 20;
        for (n20 = 0; n20 < 16; n20 = n20 + 1) 
        begin: outbit20
            assign data_11[n20 + d20*16 + c0*28*16] = data_11_array[c0][d20][n20];
        end
    endgenerate
    generate 
        localparam integer d21 = 21;
        for (n21 = 0; n21 < 16; n21 = n21 + 1) 
        begin: outbit21
            assign data_11[n21 + d21*16 + c0*28*16] = data_11_array[c0][d21][n21];
        end
    endgenerate
    generate 
        localparam integer d22 = 22;
        for (n22 = 0; n22 < 16; n22 = n22 + 1) 
        begin: outbit22
            assign data_11[n22 + d22*16 + c0*28*16] = data_11_array[c0][d22][n22];
        end
    endgenerate
    generate 
        localparam integer d23 = 23;
        for (n23 = 0; n23 < 16; n23 = n23 + 1) 
        begin: outbit23
            assign data_11[n23 + d23*16 + c0*28*16] = data_11_array[c0][d23][n23];
        end
    endgenerate
    generate 
        localparam integer d24 = 24;
        for (n24 = 0; n24 < 16; n24 = n24 + 1) 
        begin: outbit24
            assign data_11[n24 + d24*16 + c0*28*16] = data_11_array[c0][d24][n24];
        end
    endgenerate
    generate 
        localparam integer d25 = 25;
        for (n25 = 0; n25 < 16; n25 = n25 + 1) 
        begin: outbit25
            assign data_11[n25 + d25*16 + c0*28*16] = data_11_array[c0][d25][n25];
        end
    endgenerate
    generate 
        localparam integer d26 = 26;
        for (n26 = 0; n26 < 16; n26 = n26 + 1) 
        begin: outbit26
            assign data_11[n26 + d26*16 + c0*28*16] = data_11_array[c0][d26][n26];
        end
    endgenerate
    generate 
        localparam integer d27 = 27;
        for (n27 = 0; n27 < 16; n27 = n27 + 1) 
        begin: outbit27
            assign data_11[n27 + d27*16 + c0*28*16] = data_11_array[c0][d27][n27];
        end
    endgenerate
    localparam integer c1 = 1;
    generate 
        localparam integer d28 = 0;
        for (n28 = 0; n28 < 16; n28 = n28 + 1) 
        begin: outbit28
            assign data_11[n28 + d28*16 + c1*28*16] = data_11_array[c1][d28][n28];
        end
    endgenerate
    generate 
        localparam integer d29 = 1;
        for (n29 = 0; n29 < 16; n29 = n29 + 1) 
        begin: outbit29
            assign data_11[n29 + d29*16 + c1*28*16] = data_11_array[c1][d29][n29];
        end
    endgenerate
    generate 
        localparam integer d30 = 2;
        for (n30 = 0; n30 < 16; n30 = n30 + 1) 
        begin: outbit30
            assign data_11[n30 + d30*16 + c1*28*16] = data_11_array[c1][d30][n30];
        end
    endgenerate
    generate 
        localparam integer d31 = 3;
        for (n31 = 0; n31 < 16; n31 = n31 + 1) 
        begin: outbit31
            assign data_11[n31 + d31*16 + c1*28*16] = data_11_array[c1][d31][n31];
        end
    endgenerate
    generate 
        localparam integer d32 = 4;
        for (n32 = 0; n32 < 16; n32 = n32 + 1) 
        begin: outbit32
            assign data_11[n32 + d32*16 + c1*28*16] = data_11_array[c1][d32][n32];
        end
    endgenerate
    generate 
        localparam integer d33 = 5;
        for (n33 = 0; n33 < 16; n33 = n33 + 1) 
        begin: outbit33
            assign data_11[n33 + d33*16 + c1*28*16] = data_11_array[c1][d33][n33];
        end
    endgenerate
    generate 
        localparam integer d34 = 6;
        for (n34 = 0; n34 < 16; n34 = n34 + 1) 
        begin: outbit34
            assign data_11[n34 + d34*16 + c1*28*16] = data_11_array[c1][d34][n34];
        end
    endgenerate
    generate 
        localparam integer d35 = 7;
        for (n35 = 0; n35 < 16; n35 = n35 + 1) 
        begin: outbit35
            assign data_11[n35 + d35*16 + c1*28*16] = data_11_array[c1][d35][n35];
        end
    endgenerate
    generate 
        localparam integer d36 = 8;
        for (n36 = 0; n36 < 16; n36 = n36 + 1) 
        begin: outbit36
            assign data_11[n36 + d36*16 + c1*28*16] = data_11_array[c1][d36][n36];
        end
    endgenerate
    generate 
        localparam integer d37 = 9;
        for (n37 = 0; n37 < 16; n37 = n37 + 1) 
        begin: outbit37
            assign data_11[n37 + d37*16 + c1*28*16] = data_11_array[c1][d37][n37];
        end
    endgenerate
    generate 
        localparam integer d38 = 10;
        for (n38 = 0; n38 < 16; n38 = n38 + 1) 
        begin: outbit38
            assign data_11[n38 + d38*16 + c1*28*16] = data_11_array[c1][d38][n38];
        end
    endgenerate
    generate 
        localparam integer d39 = 11;
        for (n39 = 0; n39 < 16; n39 = n39 + 1) 
        begin: outbit39
            assign data_11[n39 + d39*16 + c1*28*16] = data_11_array[c1][d39][n39];
        end
    endgenerate
    generate 
        localparam integer d40 = 12;
        for (n40 = 0; n40 < 16; n40 = n40 + 1) 
        begin: outbit40
            assign data_11[n40 + d40*16 + c1*28*16] = data_11_array[c1][d40][n40];
        end
    endgenerate
    generate 
        localparam integer d41 = 13;
        for (n41 = 0; n41 < 16; n41 = n41 + 1) 
        begin: outbit41
            assign data_11[n41 + d41*16 + c1*28*16] = data_11_array[c1][d41][n41];
        end
    endgenerate
    generate 
        localparam integer d42 = 14;
        for (n42 = 0; n42 < 16; n42 = n42 + 1) 
        begin: outbit42
            assign data_11[n42 + d42*16 + c1*28*16] = data_11_array[c1][d42][n42];
        end
    endgenerate
    generate 
        localparam integer d43 = 15;
        for (n43 = 0; n43 < 16; n43 = n43 + 1) 
        begin: outbit43
            assign data_11[n43 + d43*16 + c1*28*16] = data_11_array[c1][d43][n43];
        end
    endgenerate
    generate 
        localparam integer d44 = 16;
        for (n44 = 0; n44 < 16; n44 = n44 + 1) 
        begin: outbit44
            assign data_11[n44 + d44*16 + c1*28*16] = data_11_array[c1][d44][n44];
        end
    endgenerate
    generate 
        localparam integer d45 = 17;
        for (n45 = 0; n45 < 16; n45 = n45 + 1) 
        begin: outbit45
            assign data_11[n45 + d45*16 + c1*28*16] = data_11_array[c1][d45][n45];
        end
    endgenerate
    generate 
        localparam integer d46 = 18;
        for (n46 = 0; n46 < 16; n46 = n46 + 1) 
        begin: outbit46
            assign data_11[n46 + d46*16 + c1*28*16] = data_11_array[c1][d46][n46];
        end
    endgenerate
    generate 
        localparam integer d47 = 19;
        for (n47 = 0; n47 < 16; n47 = n47 + 1) 
        begin: outbit47
            assign data_11[n47 + d47*16 + c1*28*16] = data_11_array[c1][d47][n47];
        end
    endgenerate
    generate 
        localparam integer d48 = 20;
        for (n48 = 0; n48 < 16; n48 = n48 + 1) 
        begin: outbit48
            assign data_11[n48 + d48*16 + c1*28*16] = data_11_array[c1][d48][n48];
        end
    endgenerate
    generate 
        localparam integer d49 = 21;
        for (n49 = 0; n49 < 16; n49 = n49 + 1) 
        begin: outbit49
            assign data_11[n49 + d49*16 + c1*28*16] = data_11_array[c1][d49][n49];
        end
    endgenerate
    generate 
        localparam integer d50 = 22;
        for (n50 = 0; n50 < 16; n50 = n50 + 1) 
        begin: outbit50
            assign data_11[n50 + d50*16 + c1*28*16] = data_11_array[c1][d50][n50];
        end
    endgenerate
    generate 
        localparam integer d51 = 23;
        for (n51 = 0; n51 < 16; n51 = n51 + 1) 
        begin: outbit51
            assign data_11[n51 + d51*16 + c1*28*16] = data_11_array[c1][d51][n51];
        end
    endgenerate
    generate 
        localparam integer d52 = 24;
        for (n52 = 0; n52 < 16; n52 = n52 + 1) 
        begin: outbit52
            assign data_11[n52 + d52*16 + c1*28*16] = data_11_array[c1][d52][n52];
        end
    endgenerate
    generate 
        localparam integer d53 = 25;
        for (n53 = 0; n53 < 16; n53 = n53 + 1) 
        begin: outbit53
            assign data_11[n53 + d53*16 + c1*28*16] = data_11_array[c1][d53][n53];
        end
    endgenerate
    generate 
        localparam integer d54 = 26;
        for (n54 = 0; n54 < 16; n54 = n54 + 1) 
        begin: outbit54
            assign data_11[n54 + d54*16 + c1*28*16] = data_11_array[c1][d54][n54];
        end
    endgenerate
    generate 
        localparam integer d55 = 27;
        for (n55 = 0; n55 < 16; n55 = n55 + 1) 
        begin: outbit55
            assign data_11[n55 + d55*16 + c1*28*16] = data_11_array[c1][d55][n55];
        end
    endgenerate
    localparam integer c2 = 2;
    generate 
        localparam integer d56 = 0;
        for (n56 = 0; n56 < 16; n56 = n56 + 1) 
        begin: outbit56
            assign data_11[n56 + d56*16 + c2*28*16] = data_11_array[c2][d56][n56];
        end
    endgenerate
    generate 
        localparam integer d57 = 1;
        for (n57 = 0; n57 < 16; n57 = n57 + 1) 
        begin: outbit57
            assign data_11[n57 + d57*16 + c2*28*16] = data_11_array[c2][d57][n57];
        end
    endgenerate
    generate 
        localparam integer d58 = 2;
        for (n58 = 0; n58 < 16; n58 = n58 + 1) 
        begin: outbit58
            assign data_11[n58 + d58*16 + c2*28*16] = data_11_array[c2][d58][n58];
        end
    endgenerate
    generate 
        localparam integer d59 = 3;
        for (n59 = 0; n59 < 16; n59 = n59 + 1) 
        begin: outbit59
            assign data_11[n59 + d59*16 + c2*28*16] = data_11_array[c2][d59][n59];
        end
    endgenerate
    generate 
        localparam integer d60 = 4;
        for (n60 = 0; n60 < 16; n60 = n60 + 1) 
        begin: outbit60
            assign data_11[n60 + d60*16 + c2*28*16] = data_11_array[c2][d60][n60];
        end
    endgenerate
    generate 
        localparam integer d61 = 5;
        for (n61 = 0; n61 < 16; n61 = n61 + 1) 
        begin: outbit61
            assign data_11[n61 + d61*16 + c2*28*16] = data_11_array[c2][d61][n61];
        end
    endgenerate
    generate 
        localparam integer d62 = 6;
        for (n62 = 0; n62 < 16; n62 = n62 + 1) 
        begin: outbit62
            assign data_11[n62 + d62*16 + c2*28*16] = data_11_array[c2][d62][n62];
        end
    endgenerate
    generate 
        localparam integer d63 = 7;
        for (n63 = 0; n63 < 16; n63 = n63 + 1) 
        begin: outbit63
            assign data_11[n63 + d63*16 + c2*28*16] = data_11_array[c2][d63][n63];
        end
    endgenerate
    generate 
        localparam integer d64 = 8;
        for (n64 = 0; n64 < 16; n64 = n64 + 1) 
        begin: outbit64
            assign data_11[n64 + d64*16 + c2*28*16] = data_11_array[c2][d64][n64];
        end
    endgenerate
    generate 
        localparam integer d65 = 9;
        for (n65 = 0; n65 < 16; n65 = n65 + 1) 
        begin: outbit65
            assign data_11[n65 + d65*16 + c2*28*16] = data_11_array[c2][d65][n65];
        end
    endgenerate
    generate 
        localparam integer d66 = 10;
        for (n66 = 0; n66 < 16; n66 = n66 + 1) 
        begin: outbit66
            assign data_11[n66 + d66*16 + c2*28*16] = data_11_array[c2][d66][n66];
        end
    endgenerate
    generate 
        localparam integer d67 = 11;
        for (n67 = 0; n67 < 16; n67 = n67 + 1) 
        begin: outbit67
            assign data_11[n67 + d67*16 + c2*28*16] = data_11_array[c2][d67][n67];
        end
    endgenerate
    generate 
        localparam integer d68 = 12;
        for (n68 = 0; n68 < 16; n68 = n68 + 1) 
        begin: outbit68
            assign data_11[n68 + d68*16 + c2*28*16] = data_11_array[c2][d68][n68];
        end
    endgenerate
    generate 
        localparam integer d69 = 13;
        for (n69 = 0; n69 < 16; n69 = n69 + 1) 
        begin: outbit69
            assign data_11[n69 + d69*16 + c2*28*16] = data_11_array[c2][d69][n69];
        end
    endgenerate
    generate 
        localparam integer d70 = 14;
        for (n70 = 0; n70 < 16; n70 = n70 + 1) 
        begin: outbit70
            assign data_11[n70 + d70*16 + c2*28*16] = data_11_array[c2][d70][n70];
        end
    endgenerate
    generate 
        localparam integer d71 = 15;
        for (n71 = 0; n71 < 16; n71 = n71 + 1) 
        begin: outbit71
            assign data_11[n71 + d71*16 + c2*28*16] = data_11_array[c2][d71][n71];
        end
    endgenerate
    generate 
        localparam integer d72 = 16;
        for (n72 = 0; n72 < 16; n72 = n72 + 1) 
        begin: outbit72
            assign data_11[n72 + d72*16 + c2*28*16] = data_11_array[c2][d72][n72];
        end
    endgenerate
    generate 
        localparam integer d73 = 17;
        for (n73 = 0; n73 < 16; n73 = n73 + 1) 
        begin: outbit73
            assign data_11[n73 + d73*16 + c2*28*16] = data_11_array[c2][d73][n73];
        end
    endgenerate
    generate 
        localparam integer d74 = 18;
        for (n74 = 0; n74 < 16; n74 = n74 + 1) 
        begin: outbit74
            assign data_11[n74 + d74*16 + c2*28*16] = data_11_array[c2][d74][n74];
        end
    endgenerate
    generate 
        localparam integer d75 = 19;
        for (n75 = 0; n75 < 16; n75 = n75 + 1) 
        begin: outbit75
            assign data_11[n75 + d75*16 + c2*28*16] = data_11_array[c2][d75][n75];
        end
    endgenerate
    generate 
        localparam integer d76 = 20;
        for (n76 = 0; n76 < 16; n76 = n76 + 1) 
        begin: outbit76
            assign data_11[n76 + d76*16 + c2*28*16] = data_11_array[c2][d76][n76];
        end
    endgenerate
    generate 
        localparam integer d77 = 21;
        for (n77 = 0; n77 < 16; n77 = n77 + 1) 
        begin: outbit77
            assign data_11[n77 + d77*16 + c2*28*16] = data_11_array[c2][d77][n77];
        end
    endgenerate
    generate 
        localparam integer d78 = 22;
        for (n78 = 0; n78 < 16; n78 = n78 + 1) 
        begin: outbit78
            assign data_11[n78 + d78*16 + c2*28*16] = data_11_array[c2][d78][n78];
        end
    endgenerate
    generate 
        localparam integer d79 = 23;
        for (n79 = 0; n79 < 16; n79 = n79 + 1) 
        begin: outbit79
            assign data_11[n79 + d79*16 + c2*28*16] = data_11_array[c2][d79][n79];
        end
    endgenerate
    generate 
        localparam integer d80 = 24;
        for (n80 = 0; n80 < 16; n80 = n80 + 1) 
        begin: outbit80
            assign data_11[n80 + d80*16 + c2*28*16] = data_11_array[c2][d80][n80];
        end
    endgenerate
    generate 
        localparam integer d81 = 25;
        for (n81 = 0; n81 < 16; n81 = n81 + 1) 
        begin: outbit81
            assign data_11[n81 + d81*16 + c2*28*16] = data_11_array[c2][d81][n81];
        end
    endgenerate
    generate 
        localparam integer d82 = 26;
        for (n82 = 0; n82 < 16; n82 = n82 + 1) 
        begin: outbit82
            assign data_11[n82 + d82*16 + c2*28*16] = data_11_array[c2][d82][n82];
        end
    endgenerate
    generate 
        localparam integer d83 = 27;
        for (n83 = 0; n83 < 16; n83 = n83 + 1) 
        begin: outbit83
            assign data_11[n83 + d83*16 + c2*28*16] = data_11_array[c2][d83][n83];
        end
    endgenerate
    localparam integer c3 = 3;
    generate 
        localparam integer d84 = 0;
        for (n84 = 0; n84 < 16; n84 = n84 + 1) 
        begin: outbit84
            assign data_11[n84 + d84*16 + c3*28*16] = data_11_array[c3][d84][n84];
        end
    endgenerate
    generate 
        localparam integer d85 = 1;
        for (n85 = 0; n85 < 16; n85 = n85 + 1) 
        begin: outbit85
            assign data_11[n85 + d85*16 + c3*28*16] = data_11_array[c3][d85][n85];
        end
    endgenerate
    generate 
        localparam integer d86 = 2;
        for (n86 = 0; n86 < 16; n86 = n86 + 1) 
        begin: outbit86
            assign data_11[n86 + d86*16 + c3*28*16] = data_11_array[c3][d86][n86];
        end
    endgenerate
    generate 
        localparam integer d87 = 3;
        for (n87 = 0; n87 < 16; n87 = n87 + 1) 
        begin: outbit87
            assign data_11[n87 + d87*16 + c3*28*16] = data_11_array[c3][d87][n87];
        end
    endgenerate
    generate 
        localparam integer d88 = 4;
        for (n88 = 0; n88 < 16; n88 = n88 + 1) 
        begin: outbit88
            assign data_11[n88 + d88*16 + c3*28*16] = data_11_array[c3][d88][n88];
        end
    endgenerate
    generate 
        localparam integer d89 = 5;
        for (n89 = 0; n89 < 16; n89 = n89 + 1) 
        begin: outbit89
            assign data_11[n89 + d89*16 + c3*28*16] = data_11_array[c3][d89][n89];
        end
    endgenerate
    generate 
        localparam integer d90 = 6;
        for (n90 = 0; n90 < 16; n90 = n90 + 1) 
        begin: outbit90
            assign data_11[n90 + d90*16 + c3*28*16] = data_11_array[c3][d90][n90];
        end
    endgenerate
    generate 
        localparam integer d91 = 7;
        for (n91 = 0; n91 < 16; n91 = n91 + 1) 
        begin: outbit91
            assign data_11[n91 + d91*16 + c3*28*16] = data_11_array[c3][d91][n91];
        end
    endgenerate
    generate 
        localparam integer d92 = 8;
        for (n92 = 0; n92 < 16; n92 = n92 + 1) 
        begin: outbit92
            assign data_11[n92 + d92*16 + c3*28*16] = data_11_array[c3][d92][n92];
        end
    endgenerate
    generate 
        localparam integer d93 = 9;
        for (n93 = 0; n93 < 16; n93 = n93 + 1) 
        begin: outbit93
            assign data_11[n93 + d93*16 + c3*28*16] = data_11_array[c3][d93][n93];
        end
    endgenerate
    generate 
        localparam integer d94 = 10;
        for (n94 = 0; n94 < 16; n94 = n94 + 1) 
        begin: outbit94
            assign data_11[n94 + d94*16 + c3*28*16] = data_11_array[c3][d94][n94];
        end
    endgenerate
    generate 
        localparam integer d95 = 11;
        for (n95 = 0; n95 < 16; n95 = n95 + 1) 
        begin: outbit95
            assign data_11[n95 + d95*16 + c3*28*16] = data_11_array[c3][d95][n95];
        end
    endgenerate
    generate 
        localparam integer d96 = 12;
        for (n96 = 0; n96 < 16; n96 = n96 + 1) 
        begin: outbit96
            assign data_11[n96 + d96*16 + c3*28*16] = data_11_array[c3][d96][n96];
        end
    endgenerate
    generate 
        localparam integer d97 = 13;
        for (n97 = 0; n97 < 16; n97 = n97 + 1) 
        begin: outbit97
            assign data_11[n97 + d97*16 + c3*28*16] = data_11_array[c3][d97][n97];
        end
    endgenerate
    generate 
        localparam integer d98 = 14;
        for (n98 = 0; n98 < 16; n98 = n98 + 1) 
        begin: outbit98
            assign data_11[n98 + d98*16 + c3*28*16] = data_11_array[c3][d98][n98];
        end
    endgenerate
    generate 
        localparam integer d99 = 15;
        for (n99 = 0; n99 < 16; n99 = n99 + 1) 
        begin: outbit99
            assign data_11[n99 + d99*16 + c3*28*16] = data_11_array[c3][d99][n99];
        end
    endgenerate
    generate 
        localparam integer d100 = 16;
        for (n100 = 0; n100 < 16; n100 = n100 + 1) 
        begin: outbit100
            assign data_11[n100 + d100*16 + c3*28*16] = data_11_array[c3][d100][n100];
        end
    endgenerate
    generate 
        localparam integer d101 = 17;
        for (n101 = 0; n101 < 16; n101 = n101 + 1) 
        begin: outbit101
            assign data_11[n101 + d101*16 + c3*28*16] = data_11_array[c3][d101][n101];
        end
    endgenerate
    generate 
        localparam integer d102 = 18;
        for (n102 = 0; n102 < 16; n102 = n102 + 1) 
        begin: outbit102
            assign data_11[n102 + d102*16 + c3*28*16] = data_11_array[c3][d102][n102];
        end
    endgenerate
    generate 
        localparam integer d103 = 19;
        for (n103 = 0; n103 < 16; n103 = n103 + 1) 
        begin: outbit103
            assign data_11[n103 + d103*16 + c3*28*16] = data_11_array[c3][d103][n103];
        end
    endgenerate
    generate 
        localparam integer d104 = 20;
        for (n104 = 0; n104 < 16; n104 = n104 + 1) 
        begin: outbit104
            assign data_11[n104 + d104*16 + c3*28*16] = data_11_array[c3][d104][n104];
        end
    endgenerate
    generate 
        localparam integer d105 = 21;
        for (n105 = 0; n105 < 16; n105 = n105 + 1) 
        begin: outbit105
            assign data_11[n105 + d105*16 + c3*28*16] = data_11_array[c3][d105][n105];
        end
    endgenerate
    generate 
        localparam integer d106 = 22;
        for (n106 = 0; n106 < 16; n106 = n106 + 1) 
        begin: outbit106
            assign data_11[n106 + d106*16 + c3*28*16] = data_11_array[c3][d106][n106];
        end
    endgenerate
    generate 
        localparam integer d107 = 23;
        for (n107 = 0; n107 < 16; n107 = n107 + 1) 
        begin: outbit107
            assign data_11[n107 + d107*16 + c3*28*16] = data_11_array[c3][d107][n107];
        end
    endgenerate
    generate 
        localparam integer d108 = 24;
        for (n108 = 0; n108 < 16; n108 = n108 + 1) 
        begin: outbit108
            assign data_11[n108 + d108*16 + c3*28*16] = data_11_array[c3][d108][n108];
        end
    endgenerate
    generate 
        localparam integer d109 = 25;
        for (n109 = 0; n109 < 16; n109 = n109 + 1) 
        begin: outbit109
            assign data_11[n109 + d109*16 + c3*28*16] = data_11_array[c3][d109][n109];
        end
    endgenerate
    generate 
        localparam integer d110 = 26;
        for (n110 = 0; n110 < 16; n110 = n110 + 1) 
        begin: outbit110
            assign data_11[n110 + d110*16 + c3*28*16] = data_11_array[c3][d110][n110];
        end
    endgenerate
    generate 
        localparam integer d111 = 27;
        for (n111 = 0; n111 < 16; n111 = n111 + 1) 
        begin: outbit111
            assign data_11[n111 + d111*16 + c3*28*16] = data_11_array[c3][d111][n111];
        end
    endgenerate
    localparam integer c4 = 4;
    generate 
        localparam integer d112 = 0;
        for (n112 = 0; n112 < 16; n112 = n112 + 1) 
        begin: outbit112
            assign data_11[n112 + d112*16 + c4*28*16] = data_11_array[c4][d112][n112];
        end
    endgenerate
    generate 
        localparam integer d113 = 1;
        for (n113 = 0; n113 < 16; n113 = n113 + 1) 
        begin: outbit113
            assign data_11[n113 + d113*16 + c4*28*16] = data_11_array[c4][d113][n113];
        end
    endgenerate
    generate 
        localparam integer d114 = 2;
        for (n114 = 0; n114 < 16; n114 = n114 + 1) 
        begin: outbit114
            assign data_11[n114 + d114*16 + c4*28*16] = data_11_array[c4][d114][n114];
        end
    endgenerate
    generate 
        localparam integer d115 = 3;
        for (n115 = 0; n115 < 16; n115 = n115 + 1) 
        begin: outbit115
            assign data_11[n115 + d115*16 + c4*28*16] = data_11_array[c4][d115][n115];
        end
    endgenerate
    generate 
        localparam integer d116 = 4;
        for (n116 = 0; n116 < 16; n116 = n116 + 1) 
        begin: outbit116
            assign data_11[n116 + d116*16 + c4*28*16] = data_11_array[c4][d116][n116];
        end
    endgenerate
    generate 
        localparam integer d117 = 5;
        for (n117 = 0; n117 < 16; n117 = n117 + 1) 
        begin: outbit117
            assign data_11[n117 + d117*16 + c4*28*16] = data_11_array[c4][d117][n117];
        end
    endgenerate
    generate 
        localparam integer d118 = 6;
        for (n118 = 0; n118 < 16; n118 = n118 + 1) 
        begin: outbit118
            assign data_11[n118 + d118*16 + c4*28*16] = data_11_array[c4][d118][n118];
        end
    endgenerate
    generate 
        localparam integer d119 = 7;
        for (n119 = 0; n119 < 16; n119 = n119 + 1) 
        begin: outbit119
            assign data_11[n119 + d119*16 + c4*28*16] = data_11_array[c4][d119][n119];
        end
    endgenerate
    generate 
        localparam integer d120 = 8;
        for (n120 = 0; n120 < 16; n120 = n120 + 1) 
        begin: outbit120
            assign data_11[n120 + d120*16 + c4*28*16] = data_11_array[c4][d120][n120];
        end
    endgenerate
    generate 
        localparam integer d121 = 9;
        for (n121 = 0; n121 < 16; n121 = n121 + 1) 
        begin: outbit121
            assign data_11[n121 + d121*16 + c4*28*16] = data_11_array[c4][d121][n121];
        end
    endgenerate
    generate 
        localparam integer d122 = 10;
        for (n122 = 0; n122 < 16; n122 = n122 + 1) 
        begin: outbit122
            assign data_11[n122 + d122*16 + c4*28*16] = data_11_array[c4][d122][n122];
        end
    endgenerate
    generate 
        localparam integer d123 = 11;
        for (n123 = 0; n123 < 16; n123 = n123 + 1) 
        begin: outbit123
            assign data_11[n123 + d123*16 + c4*28*16] = data_11_array[c4][d123][n123];
        end
    endgenerate
    generate 
        localparam integer d124 = 12;
        for (n124 = 0; n124 < 16; n124 = n124 + 1) 
        begin: outbit124
            assign data_11[n124 + d124*16 + c4*28*16] = data_11_array[c4][d124][n124];
        end
    endgenerate
    generate 
        localparam integer d125 = 13;
        for (n125 = 0; n125 < 16; n125 = n125 + 1) 
        begin: outbit125
            assign data_11[n125 + d125*16 + c4*28*16] = data_11_array[c4][d125][n125];
        end
    endgenerate
    generate 
        localparam integer d126 = 14;
        for (n126 = 0; n126 < 16; n126 = n126 + 1) 
        begin: outbit126
            assign data_11[n126 + d126*16 + c4*28*16] = data_11_array[c4][d126][n126];
        end
    endgenerate
    generate 
        localparam integer d127 = 15;
        for (n127 = 0; n127 < 16; n127 = n127 + 1) 
        begin: outbit127
            assign data_11[n127 + d127*16 + c4*28*16] = data_11_array[c4][d127][n127];
        end
    endgenerate
    generate 
        localparam integer d128 = 16;
        for (n128 = 0; n128 < 16; n128 = n128 + 1) 
        begin: outbit128
            assign data_11[n128 + d128*16 + c4*28*16] = data_11_array[c4][d128][n128];
        end
    endgenerate
    generate 
        localparam integer d129 = 17;
        for (n129 = 0; n129 < 16; n129 = n129 + 1) 
        begin: outbit129
            assign data_11[n129 + d129*16 + c4*28*16] = data_11_array[c4][d129][n129];
        end
    endgenerate
    generate 
        localparam integer d130 = 18;
        for (n130 = 0; n130 < 16; n130 = n130 + 1) 
        begin: outbit130
            assign data_11[n130 + d130*16 + c4*28*16] = data_11_array[c4][d130][n130];
        end
    endgenerate
    generate 
        localparam integer d131 = 19;
        for (n131 = 0; n131 < 16; n131 = n131 + 1) 
        begin: outbit131
            assign data_11[n131 + d131*16 + c4*28*16] = data_11_array[c4][d131][n131];
        end
    endgenerate
    generate 
        localparam integer d132 = 20;
        for (n132 = 0; n132 < 16; n132 = n132 + 1) 
        begin: outbit132
            assign data_11[n132 + d132*16 + c4*28*16] = data_11_array[c4][d132][n132];
        end
    endgenerate
    generate 
        localparam integer d133 = 21;
        for (n133 = 0; n133 < 16; n133 = n133 + 1) 
        begin: outbit133
            assign data_11[n133 + d133*16 + c4*28*16] = data_11_array[c4][d133][n133];
        end
    endgenerate
    generate 
        localparam integer d134 = 22;
        for (n134 = 0; n134 < 16; n134 = n134 + 1) 
        begin: outbit134
            assign data_11[n134 + d134*16 + c4*28*16] = data_11_array[c4][d134][n134];
        end
    endgenerate
    generate 
        localparam integer d135 = 23;
        for (n135 = 0; n135 < 16; n135 = n135 + 1) 
        begin: outbit135
            assign data_11[n135 + d135*16 + c4*28*16] = data_11_array[c4][d135][n135];
        end
    endgenerate
    generate 
        localparam integer d136 = 24;
        for (n136 = 0; n136 < 16; n136 = n136 + 1) 
        begin: outbit136
            assign data_11[n136 + d136*16 + c4*28*16] = data_11_array[c4][d136][n136];
        end
    endgenerate
    generate 
        localparam integer d137 = 25;
        for (n137 = 0; n137 < 16; n137 = n137 + 1) 
        begin: outbit137
            assign data_11[n137 + d137*16 + c4*28*16] = data_11_array[c4][d137][n137];
        end
    endgenerate
    generate 
        localparam integer d138 = 26;
        for (n138 = 0; n138 < 16; n138 = n138 + 1) 
        begin: outbit138
            assign data_11[n138 + d138*16 + c4*28*16] = data_11_array[c4][d138][n138];
        end
    endgenerate
    generate 
        localparam integer d139 = 27;
        for (n139 = 0; n139 < 16; n139 = n139 + 1) 
        begin: outbit139
            assign data_11[n139 + d139*16 + c4*28*16] = data_11_array[c4][d139][n139];
        end
    endgenerate
    localparam integer c5 = 5;
    generate 
        localparam integer d140 = 0;
        for (n140 = 0; n140 < 16; n140 = n140 + 1) 
        begin: outbit140
            assign data_11[n140 + d140*16 + c5*28*16] = data_11_array[c5][d140][n140];
        end
    endgenerate
    generate 
        localparam integer d141 = 1;
        for (n141 = 0; n141 < 16; n141 = n141 + 1) 
        begin: outbit141
            assign data_11[n141 + d141*16 + c5*28*16] = data_11_array[c5][d141][n141];
        end
    endgenerate
    generate 
        localparam integer d142 = 2;
        for (n142 = 0; n142 < 16; n142 = n142 + 1) 
        begin: outbit142
            assign data_11[n142 + d142*16 + c5*28*16] = data_11_array[c5][d142][n142];
        end
    endgenerate
    generate 
        localparam integer d143 = 3;
        for (n143 = 0; n143 < 16; n143 = n143 + 1) 
        begin: outbit143
            assign data_11[n143 + d143*16 + c5*28*16] = data_11_array[c5][d143][n143];
        end
    endgenerate
    generate 
        localparam integer d144 = 4;
        for (n144 = 0; n144 < 16; n144 = n144 + 1) 
        begin: outbit144
            assign data_11[n144 + d144*16 + c5*28*16] = data_11_array[c5][d144][n144];
        end
    endgenerate
    generate 
        localparam integer d145 = 5;
        for (n145 = 0; n145 < 16; n145 = n145 + 1) 
        begin: outbit145
            assign data_11[n145 + d145*16 + c5*28*16] = data_11_array[c5][d145][n145];
        end
    endgenerate
    generate 
        localparam integer d146 = 6;
        for (n146 = 0; n146 < 16; n146 = n146 + 1) 
        begin: outbit146
            assign data_11[n146 + d146*16 + c5*28*16] = data_11_array[c5][d146][n146];
        end
    endgenerate
    generate 
        localparam integer d147 = 7;
        for (n147 = 0; n147 < 16; n147 = n147 + 1) 
        begin: outbit147
            assign data_11[n147 + d147*16 + c5*28*16] = data_11_array[c5][d147][n147];
        end
    endgenerate
    generate 
        localparam integer d148 = 8;
        for (n148 = 0; n148 < 16; n148 = n148 + 1) 
        begin: outbit148
            assign data_11[n148 + d148*16 + c5*28*16] = data_11_array[c5][d148][n148];
        end
    endgenerate
    generate 
        localparam integer d149 = 9;
        for (n149 = 0; n149 < 16; n149 = n149 + 1) 
        begin: outbit149
            assign data_11[n149 + d149*16 + c5*28*16] = data_11_array[c5][d149][n149];
        end
    endgenerate
    generate 
        localparam integer d150 = 10;
        for (n150 = 0; n150 < 16; n150 = n150 + 1) 
        begin: outbit150
            assign data_11[n150 + d150*16 + c5*28*16] = data_11_array[c5][d150][n150];
        end
    endgenerate
    generate 
        localparam integer d151 = 11;
        for (n151 = 0; n151 < 16; n151 = n151 + 1) 
        begin: outbit151
            assign data_11[n151 + d151*16 + c5*28*16] = data_11_array[c5][d151][n151];
        end
    endgenerate
    generate 
        localparam integer d152 = 12;
        for (n152 = 0; n152 < 16; n152 = n152 + 1) 
        begin: outbit152
            assign data_11[n152 + d152*16 + c5*28*16] = data_11_array[c5][d152][n152];
        end
    endgenerate
    generate 
        localparam integer d153 = 13;
        for (n153 = 0; n153 < 16; n153 = n153 + 1) 
        begin: outbit153
            assign data_11[n153 + d153*16 + c5*28*16] = data_11_array[c5][d153][n153];
        end
    endgenerate
    generate 
        localparam integer d154 = 14;
        for (n154 = 0; n154 < 16; n154 = n154 + 1) 
        begin: outbit154
            assign data_11[n154 + d154*16 + c5*28*16] = data_11_array[c5][d154][n154];
        end
    endgenerate
    generate 
        localparam integer d155 = 15;
        for (n155 = 0; n155 < 16; n155 = n155 + 1) 
        begin: outbit155
            assign data_11[n155 + d155*16 + c5*28*16] = data_11_array[c5][d155][n155];
        end
    endgenerate
    generate 
        localparam integer d156 = 16;
        for (n156 = 0; n156 < 16; n156 = n156 + 1) 
        begin: outbit156
            assign data_11[n156 + d156*16 + c5*28*16] = data_11_array[c5][d156][n156];
        end
    endgenerate
    generate 
        localparam integer d157 = 17;
        for (n157 = 0; n157 < 16; n157 = n157 + 1) 
        begin: outbit157
            assign data_11[n157 + d157*16 + c5*28*16] = data_11_array[c5][d157][n157];
        end
    endgenerate
    generate 
        localparam integer d158 = 18;
        for (n158 = 0; n158 < 16; n158 = n158 + 1) 
        begin: outbit158
            assign data_11[n158 + d158*16 + c5*28*16] = data_11_array[c5][d158][n158];
        end
    endgenerate
    generate 
        localparam integer d159 = 19;
        for (n159 = 0; n159 < 16; n159 = n159 + 1) 
        begin: outbit159
            assign data_11[n159 + d159*16 + c5*28*16] = data_11_array[c5][d159][n159];
        end
    endgenerate
    generate 
        localparam integer d160 = 20;
        for (n160 = 0; n160 < 16; n160 = n160 + 1) 
        begin: outbit160
            assign data_11[n160 + d160*16 + c5*28*16] = data_11_array[c5][d160][n160];
        end
    endgenerate
    generate 
        localparam integer d161 = 21;
        for (n161 = 0; n161 < 16; n161 = n161 + 1) 
        begin: outbit161
            assign data_11[n161 + d161*16 + c5*28*16] = data_11_array[c5][d161][n161];
        end
    endgenerate
    generate 
        localparam integer d162 = 22;
        for (n162 = 0; n162 < 16; n162 = n162 + 1) 
        begin: outbit162
            assign data_11[n162 + d162*16 + c5*28*16] = data_11_array[c5][d162][n162];
        end
    endgenerate
    generate 
        localparam integer d163 = 23;
        for (n163 = 0; n163 < 16; n163 = n163 + 1) 
        begin: outbit163
            assign data_11[n163 + d163*16 + c5*28*16] = data_11_array[c5][d163][n163];
        end
    endgenerate
    generate 
        localparam integer d164 = 24;
        for (n164 = 0; n164 < 16; n164 = n164 + 1) 
        begin: outbit164
            assign data_11[n164 + d164*16 + c5*28*16] = data_11_array[c5][d164][n164];
        end
    endgenerate
    generate 
        localparam integer d165 = 25;
        for (n165 = 0; n165 < 16; n165 = n165 + 1) 
        begin: outbit165
            assign data_11[n165 + d165*16 + c5*28*16] = data_11_array[c5][d165][n165];
        end
    endgenerate
    generate 
        localparam integer d166 = 26;
        for (n166 = 0; n166 < 16; n166 = n166 + 1) 
        begin: outbit166
            assign data_11[n166 + d166*16 + c5*28*16] = data_11_array[c5][d166][n166];
        end
    endgenerate
    generate 
        localparam integer d167 = 27;
        for (n167 = 0; n167 < 16; n167 = n167 + 1) 
        begin: outbit167
            assign data_11[n167 + d167*16 + c5*28*16] = data_11_array[c5][d167][n167];
        end
    endgenerate
    localparam integer c6 = 6;
    generate 
        localparam integer d168 = 0;
        for (n168 = 0; n168 < 16; n168 = n168 + 1) 
        begin: outbit168
            assign data_11[n168 + d168*16 + c6*28*16] = data_11_array[c6][d168][n168];
        end
    endgenerate
    generate 
        localparam integer d169 = 1;
        for (n169 = 0; n169 < 16; n169 = n169 + 1) 
        begin: outbit169
            assign data_11[n169 + d169*16 + c6*28*16] = data_11_array[c6][d169][n169];
        end
    endgenerate
    generate 
        localparam integer d170 = 2;
        for (n170 = 0; n170 < 16; n170 = n170 + 1) 
        begin: outbit170
            assign data_11[n170 + d170*16 + c6*28*16] = data_11_array[c6][d170][n170];
        end
    endgenerate
    generate 
        localparam integer d171 = 3;
        for (n171 = 0; n171 < 16; n171 = n171 + 1) 
        begin: outbit171
            assign data_11[n171 + d171*16 + c6*28*16] = data_11_array[c6][d171][n171];
        end
    endgenerate
    generate 
        localparam integer d172 = 4;
        for (n172 = 0; n172 < 16; n172 = n172 + 1) 
        begin: outbit172
            assign data_11[n172 + d172*16 + c6*28*16] = data_11_array[c6][d172][n172];
        end
    endgenerate
    generate 
        localparam integer d173 = 5;
        for (n173 = 0; n173 < 16; n173 = n173 + 1) 
        begin: outbit173
            assign data_11[n173 + d173*16 + c6*28*16] = data_11_array[c6][d173][n173];
        end
    endgenerate
    generate 
        localparam integer d174 = 6;
        for (n174 = 0; n174 < 16; n174 = n174 + 1) 
        begin: outbit174
            assign data_11[n174 + d174*16 + c6*28*16] = data_11_array[c6][d174][n174];
        end
    endgenerate
    generate 
        localparam integer d175 = 7;
        for (n175 = 0; n175 < 16; n175 = n175 + 1) 
        begin: outbit175
            assign data_11[n175 + d175*16 + c6*28*16] = data_11_array[c6][d175][n175];
        end
    endgenerate
    generate 
        localparam integer d176 = 8;
        for (n176 = 0; n176 < 16; n176 = n176 + 1) 
        begin: outbit176
            assign data_11[n176 + d176*16 + c6*28*16] = data_11_array[c6][d176][n176];
        end
    endgenerate
    generate 
        localparam integer d177 = 9;
        for (n177 = 0; n177 < 16; n177 = n177 + 1) 
        begin: outbit177
            assign data_11[n177 + d177*16 + c6*28*16] = data_11_array[c6][d177][n177];
        end
    endgenerate
    generate 
        localparam integer d178 = 10;
        for (n178 = 0; n178 < 16; n178 = n178 + 1) 
        begin: outbit178
            assign data_11[n178 + d178*16 + c6*28*16] = data_11_array[c6][d178][n178];
        end
    endgenerate
    generate 
        localparam integer d179 = 11;
        for (n179 = 0; n179 < 16; n179 = n179 + 1) 
        begin: outbit179
            assign data_11[n179 + d179*16 + c6*28*16] = data_11_array[c6][d179][n179];
        end
    endgenerate
    generate 
        localparam integer d180 = 12;
        for (n180 = 0; n180 < 16; n180 = n180 + 1) 
        begin: outbit180
            assign data_11[n180 + d180*16 + c6*28*16] = data_11_array[c6][d180][n180];
        end
    endgenerate
    generate 
        localparam integer d181 = 13;
        for (n181 = 0; n181 < 16; n181 = n181 + 1) 
        begin: outbit181
            assign data_11[n181 + d181*16 + c6*28*16] = data_11_array[c6][d181][n181];
        end
    endgenerate
    generate 
        localparam integer d182 = 14;
        for (n182 = 0; n182 < 16; n182 = n182 + 1) 
        begin: outbit182
            assign data_11[n182 + d182*16 + c6*28*16] = data_11_array[c6][d182][n182];
        end
    endgenerate
    generate 
        localparam integer d183 = 15;
        for (n183 = 0; n183 < 16; n183 = n183 + 1) 
        begin: outbit183
            assign data_11[n183 + d183*16 + c6*28*16] = data_11_array[c6][d183][n183];
        end
    endgenerate
    generate 
        localparam integer d184 = 16;
        for (n184 = 0; n184 < 16; n184 = n184 + 1) 
        begin: outbit184
            assign data_11[n184 + d184*16 + c6*28*16] = data_11_array[c6][d184][n184];
        end
    endgenerate
    generate 
        localparam integer d185 = 17;
        for (n185 = 0; n185 < 16; n185 = n185 + 1) 
        begin: outbit185
            assign data_11[n185 + d185*16 + c6*28*16] = data_11_array[c6][d185][n185];
        end
    endgenerate
    generate 
        localparam integer d186 = 18;
        for (n186 = 0; n186 < 16; n186 = n186 + 1) 
        begin: outbit186
            assign data_11[n186 + d186*16 + c6*28*16] = data_11_array[c6][d186][n186];
        end
    endgenerate
    generate 
        localparam integer d187 = 19;
        for (n187 = 0; n187 < 16; n187 = n187 + 1) 
        begin: outbit187
            assign data_11[n187 + d187*16 + c6*28*16] = data_11_array[c6][d187][n187];
        end
    endgenerate
    generate 
        localparam integer d188 = 20;
        for (n188 = 0; n188 < 16; n188 = n188 + 1) 
        begin: outbit188
            assign data_11[n188 + d188*16 + c6*28*16] = data_11_array[c6][d188][n188];
        end
    endgenerate
    generate 
        localparam integer d189 = 21;
        for (n189 = 0; n189 < 16; n189 = n189 + 1) 
        begin: outbit189
            assign data_11[n189 + d189*16 + c6*28*16] = data_11_array[c6][d189][n189];
        end
    endgenerate
    generate 
        localparam integer d190 = 22;
        for (n190 = 0; n190 < 16; n190 = n190 + 1) 
        begin: outbit190
            assign data_11[n190 + d190*16 + c6*28*16] = data_11_array[c6][d190][n190];
        end
    endgenerate
    generate 
        localparam integer d191 = 23;
        for (n191 = 0; n191 < 16; n191 = n191 + 1) 
        begin: outbit191
            assign data_11[n191 + d191*16 + c6*28*16] = data_11_array[c6][d191][n191];
        end
    endgenerate
    generate 
        localparam integer d192 = 24;
        for (n192 = 0; n192 < 16; n192 = n192 + 1) 
        begin: outbit192
            assign data_11[n192 + d192*16 + c6*28*16] = data_11_array[c6][d192][n192];
        end
    endgenerate
    generate 
        localparam integer d193 = 25;
        for (n193 = 0; n193 < 16; n193 = n193 + 1) 
        begin: outbit193
            assign data_11[n193 + d193*16 + c6*28*16] = data_11_array[c6][d193][n193];
        end
    endgenerate
    generate 
        localparam integer d194 = 26;
        for (n194 = 0; n194 < 16; n194 = n194 + 1) 
        begin: outbit194
            assign data_11[n194 + d194*16 + c6*28*16] = data_11_array[c6][d194][n194];
        end
    endgenerate
    generate 
        localparam integer d195 = 27;
        for (n195 = 0; n195 < 16; n195 = n195 + 1) 
        begin: outbit195
            assign data_11[n195 + d195*16 + c6*28*16] = data_11_array[c6][d195][n195];
        end
    endgenerate
    localparam integer c7 = 7;
    generate 
        localparam integer d196 = 0;
        for (n196 = 0; n196 < 16; n196 = n196 + 1) 
        begin: outbit196
            assign data_11[n196 + d196*16 + c7*28*16] = data_11_array[c7][d196][n196];
        end
    endgenerate
    generate 
        localparam integer d197 = 1;
        for (n197 = 0; n197 < 16; n197 = n197 + 1) 
        begin: outbit197
            assign data_11[n197 + d197*16 + c7*28*16] = data_11_array[c7][d197][n197];
        end
    endgenerate
    generate 
        localparam integer d198 = 2;
        for (n198 = 0; n198 < 16; n198 = n198 + 1) 
        begin: outbit198
            assign data_11[n198 + d198*16 + c7*28*16] = data_11_array[c7][d198][n198];
        end
    endgenerate
    generate 
        localparam integer d199 = 3;
        for (n199 = 0; n199 < 16; n199 = n199 + 1) 
        begin: outbit199
            assign data_11[n199 + d199*16 + c7*28*16] = data_11_array[c7][d199][n199];
        end
    endgenerate
    generate 
        localparam integer d200 = 4;
        for (n200 = 0; n200 < 16; n200 = n200 + 1) 
        begin: outbit200
            assign data_11[n200 + d200*16 + c7*28*16] = data_11_array[c7][d200][n200];
        end
    endgenerate
    generate 
        localparam integer d201 = 5;
        for (n201 = 0; n201 < 16; n201 = n201 + 1) 
        begin: outbit201
            assign data_11[n201 + d201*16 + c7*28*16] = data_11_array[c7][d201][n201];
        end
    endgenerate
    generate 
        localparam integer d202 = 6;
        for (n202 = 0; n202 < 16; n202 = n202 + 1) 
        begin: outbit202
            assign data_11[n202 + d202*16 + c7*28*16] = data_11_array[c7][d202][n202];
        end
    endgenerate
    generate 
        localparam integer d203 = 7;
        for (n203 = 0; n203 < 16; n203 = n203 + 1) 
        begin: outbit203
            assign data_11[n203 + d203*16 + c7*28*16] = data_11_array[c7][d203][n203];
        end
    endgenerate
    generate 
        localparam integer d204 = 8;
        for (n204 = 0; n204 < 16; n204 = n204 + 1) 
        begin: outbit204
            assign data_11[n204 + d204*16 + c7*28*16] = data_11_array[c7][d204][n204];
        end
    endgenerate
    generate 
        localparam integer d205 = 9;
        for (n205 = 0; n205 < 16; n205 = n205 + 1) 
        begin: outbit205
            assign data_11[n205 + d205*16 + c7*28*16] = data_11_array[c7][d205][n205];
        end
    endgenerate
    generate 
        localparam integer d206 = 10;
        for (n206 = 0; n206 < 16; n206 = n206 + 1) 
        begin: outbit206
            assign data_11[n206 + d206*16 + c7*28*16] = data_11_array[c7][d206][n206];
        end
    endgenerate
    generate 
        localparam integer d207 = 11;
        for (n207 = 0; n207 < 16; n207 = n207 + 1) 
        begin: outbit207
            assign data_11[n207 + d207*16 + c7*28*16] = data_11_array[c7][d207][n207];
        end
    endgenerate
    generate 
        localparam integer d208 = 12;
        for (n208 = 0; n208 < 16; n208 = n208 + 1) 
        begin: outbit208
            assign data_11[n208 + d208*16 + c7*28*16] = data_11_array[c7][d208][n208];
        end
    endgenerate
    generate 
        localparam integer d209 = 13;
        for (n209 = 0; n209 < 16; n209 = n209 + 1) 
        begin: outbit209
            assign data_11[n209 + d209*16 + c7*28*16] = data_11_array[c7][d209][n209];
        end
    endgenerate
    generate 
        localparam integer d210 = 14;
        for (n210 = 0; n210 < 16; n210 = n210 + 1) 
        begin: outbit210
            assign data_11[n210 + d210*16 + c7*28*16] = data_11_array[c7][d210][n210];
        end
    endgenerate
    generate 
        localparam integer d211 = 15;
        for (n211 = 0; n211 < 16; n211 = n211 + 1) 
        begin: outbit211
            assign data_11[n211 + d211*16 + c7*28*16] = data_11_array[c7][d211][n211];
        end
    endgenerate
    generate 
        localparam integer d212 = 16;
        for (n212 = 0; n212 < 16; n212 = n212 + 1) 
        begin: outbit212
            assign data_11[n212 + d212*16 + c7*28*16] = data_11_array[c7][d212][n212];
        end
    endgenerate
    generate 
        localparam integer d213 = 17;
        for (n213 = 0; n213 < 16; n213 = n213 + 1) 
        begin: outbit213
            assign data_11[n213 + d213*16 + c7*28*16] = data_11_array[c7][d213][n213];
        end
    endgenerate
    generate 
        localparam integer d214 = 18;
        for (n214 = 0; n214 < 16; n214 = n214 + 1) 
        begin: outbit214
            assign data_11[n214 + d214*16 + c7*28*16] = data_11_array[c7][d214][n214];
        end
    endgenerate
    generate 
        localparam integer d215 = 19;
        for (n215 = 0; n215 < 16; n215 = n215 + 1) 
        begin: outbit215
            assign data_11[n215 + d215*16 + c7*28*16] = data_11_array[c7][d215][n215];
        end
    endgenerate
    generate 
        localparam integer d216 = 20;
        for (n216 = 0; n216 < 16; n216 = n216 + 1) 
        begin: outbit216
            assign data_11[n216 + d216*16 + c7*28*16] = data_11_array[c7][d216][n216];
        end
    endgenerate
    generate 
        localparam integer d217 = 21;
        for (n217 = 0; n217 < 16; n217 = n217 + 1) 
        begin: outbit217
            assign data_11[n217 + d217*16 + c7*28*16] = data_11_array[c7][d217][n217];
        end
    endgenerate
    generate 
        localparam integer d218 = 22;
        for (n218 = 0; n218 < 16; n218 = n218 + 1) 
        begin: outbit218
            assign data_11[n218 + d218*16 + c7*28*16] = data_11_array[c7][d218][n218];
        end
    endgenerate
    generate 
        localparam integer d219 = 23;
        for (n219 = 0; n219 < 16; n219 = n219 + 1) 
        begin: outbit219
            assign data_11[n219 + d219*16 + c7*28*16] = data_11_array[c7][d219][n219];
        end
    endgenerate
    generate 
        localparam integer d220 = 24;
        for (n220 = 0; n220 < 16; n220 = n220 + 1) 
        begin: outbit220
            assign data_11[n220 + d220*16 + c7*28*16] = data_11_array[c7][d220][n220];
        end
    endgenerate
    generate 
        localparam integer d221 = 25;
        for (n221 = 0; n221 < 16; n221 = n221 + 1) 
        begin: outbit221
            assign data_11[n221 + d221*16 + c7*28*16] = data_11_array[c7][d221][n221];
        end
    endgenerate
    generate 
        localparam integer d222 = 26;
        for (n222 = 0; n222 < 16; n222 = n222 + 1) 
        begin: outbit222
            assign data_11[n222 + d222*16 + c7*28*16] = data_11_array[c7][d222][n222];
        end
    endgenerate
    generate 
        localparam integer d223 = 27;
        for (n223 = 0; n223 < 16; n223 = n223 + 1) 
        begin: outbit223
            assign data_11[n223 + d223*16 + c7*28*16] = data_11_array[c7][d223][n223];
        end
    endgenerate
    localparam integer c8 = 8;
    generate 
        localparam integer d224 = 0;
        for (n224 = 0; n224 < 16; n224 = n224 + 1) 
        begin: outbit224
            assign data_11[n224 + d224*16 + c8*28*16] = data_11_array[c8][d224][n224];
        end
    endgenerate
    generate 
        localparam integer d225 = 1;
        for (n225 = 0; n225 < 16; n225 = n225 + 1) 
        begin: outbit225
            assign data_11[n225 + d225*16 + c8*28*16] = data_11_array[c8][d225][n225];
        end
    endgenerate
    generate 
        localparam integer d226 = 2;
        for (n226 = 0; n226 < 16; n226 = n226 + 1) 
        begin: outbit226
            assign data_11[n226 + d226*16 + c8*28*16] = data_11_array[c8][d226][n226];
        end
    endgenerate
    generate 
        localparam integer d227 = 3;
        for (n227 = 0; n227 < 16; n227 = n227 + 1) 
        begin: outbit227
            assign data_11[n227 + d227*16 + c8*28*16] = data_11_array[c8][d227][n227];
        end
    endgenerate
    generate 
        localparam integer d228 = 4;
        for (n228 = 0; n228 < 16; n228 = n228 + 1) 
        begin: outbit228
            assign data_11[n228 + d228*16 + c8*28*16] = data_11_array[c8][d228][n228];
        end
    endgenerate
    generate 
        localparam integer d229 = 5;
        for (n229 = 0; n229 < 16; n229 = n229 + 1) 
        begin: outbit229
            assign data_11[n229 + d229*16 + c8*28*16] = data_11_array[c8][d229][n229];
        end
    endgenerate
    generate 
        localparam integer d230 = 6;
        for (n230 = 0; n230 < 16; n230 = n230 + 1) 
        begin: outbit230
            assign data_11[n230 + d230*16 + c8*28*16] = data_11_array[c8][d230][n230];
        end
    endgenerate
    generate 
        localparam integer d231 = 7;
        for (n231 = 0; n231 < 16; n231 = n231 + 1) 
        begin: outbit231
            assign data_11[n231 + d231*16 + c8*28*16] = data_11_array[c8][d231][n231];
        end
    endgenerate
    generate 
        localparam integer d232 = 8;
        for (n232 = 0; n232 < 16; n232 = n232 + 1) 
        begin: outbit232
            assign data_11[n232 + d232*16 + c8*28*16] = data_11_array[c8][d232][n232];
        end
    endgenerate
    generate 
        localparam integer d233 = 9;
        for (n233 = 0; n233 < 16; n233 = n233 + 1) 
        begin: outbit233
            assign data_11[n233 + d233*16 + c8*28*16] = data_11_array[c8][d233][n233];
        end
    endgenerate
    generate 
        localparam integer d234 = 10;
        for (n234 = 0; n234 < 16; n234 = n234 + 1) 
        begin: outbit234
            assign data_11[n234 + d234*16 + c8*28*16] = data_11_array[c8][d234][n234];
        end
    endgenerate
    generate 
        localparam integer d235 = 11;
        for (n235 = 0; n235 < 16; n235 = n235 + 1) 
        begin: outbit235
            assign data_11[n235 + d235*16 + c8*28*16] = data_11_array[c8][d235][n235];
        end
    endgenerate
    generate 
        localparam integer d236 = 12;
        for (n236 = 0; n236 < 16; n236 = n236 + 1) 
        begin: outbit236
            assign data_11[n236 + d236*16 + c8*28*16] = data_11_array[c8][d236][n236];
        end
    endgenerate
    generate 
        localparam integer d237 = 13;
        for (n237 = 0; n237 < 16; n237 = n237 + 1) 
        begin: outbit237
            assign data_11[n237 + d237*16 + c8*28*16] = data_11_array[c8][d237][n237];
        end
    endgenerate
    generate 
        localparam integer d238 = 14;
        for (n238 = 0; n238 < 16; n238 = n238 + 1) 
        begin: outbit238
            assign data_11[n238 + d238*16 + c8*28*16] = data_11_array[c8][d238][n238];
        end
    endgenerate
    generate 
        localparam integer d239 = 15;
        for (n239 = 0; n239 < 16; n239 = n239 + 1) 
        begin: outbit239
            assign data_11[n239 + d239*16 + c8*28*16] = data_11_array[c8][d239][n239];
        end
    endgenerate
    generate 
        localparam integer d240 = 16;
        for (n240 = 0; n240 < 16; n240 = n240 + 1) 
        begin: outbit240
            assign data_11[n240 + d240*16 + c8*28*16] = data_11_array[c8][d240][n240];
        end
    endgenerate
    generate 
        localparam integer d241 = 17;
        for (n241 = 0; n241 < 16; n241 = n241 + 1) 
        begin: outbit241
            assign data_11[n241 + d241*16 + c8*28*16] = data_11_array[c8][d241][n241];
        end
    endgenerate
    generate 
        localparam integer d242 = 18;
        for (n242 = 0; n242 < 16; n242 = n242 + 1) 
        begin: outbit242
            assign data_11[n242 + d242*16 + c8*28*16] = data_11_array[c8][d242][n242];
        end
    endgenerate
    generate 
        localparam integer d243 = 19;
        for (n243 = 0; n243 < 16; n243 = n243 + 1) 
        begin: outbit243
            assign data_11[n243 + d243*16 + c8*28*16] = data_11_array[c8][d243][n243];
        end
    endgenerate
    generate 
        localparam integer d244 = 20;
        for (n244 = 0; n244 < 16; n244 = n244 + 1) 
        begin: outbit244
            assign data_11[n244 + d244*16 + c8*28*16] = data_11_array[c8][d244][n244];
        end
    endgenerate
    generate 
        localparam integer d245 = 21;
        for (n245 = 0; n245 < 16; n245 = n245 + 1) 
        begin: outbit245
            assign data_11[n245 + d245*16 + c8*28*16] = data_11_array[c8][d245][n245];
        end
    endgenerate
    generate 
        localparam integer d246 = 22;
        for (n246 = 0; n246 < 16; n246 = n246 + 1) 
        begin: outbit246
            assign data_11[n246 + d246*16 + c8*28*16] = data_11_array[c8][d246][n246];
        end
    endgenerate
    generate 
        localparam integer d247 = 23;
        for (n247 = 0; n247 < 16; n247 = n247 + 1) 
        begin: outbit247
            assign data_11[n247 + d247*16 + c8*28*16] = data_11_array[c8][d247][n247];
        end
    endgenerate
    generate 
        localparam integer d248 = 24;
        for (n248 = 0; n248 < 16; n248 = n248 + 1) 
        begin: outbit248
            assign data_11[n248 + d248*16 + c8*28*16] = data_11_array[c8][d248][n248];
        end
    endgenerate
    generate 
        localparam integer d249 = 25;
        for (n249 = 0; n249 < 16; n249 = n249 + 1) 
        begin: outbit249
            assign data_11[n249 + d249*16 + c8*28*16] = data_11_array[c8][d249][n249];
        end
    endgenerate
    generate 
        localparam integer d250 = 26;
        for (n250 = 0; n250 < 16; n250 = n250 + 1) 
        begin: outbit250
            assign data_11[n250 + d250*16 + c8*28*16] = data_11_array[c8][d250][n250];
        end
    endgenerate
    generate 
        localparam integer d251 = 27;
        for (n251 = 0; n251 < 16; n251 = n251 + 1) 
        begin: outbit251
            assign data_11[n251 + d251*16 + c8*28*16] = data_11_array[c8][d251][n251];
        end
    endgenerate
    localparam integer c9 = 9;
    generate 
        localparam integer d252 = 0;
        for (n252 = 0; n252 < 16; n252 = n252 + 1) 
        begin: outbit252
            assign data_11[n252 + d252*16 + c9*28*16] = data_11_array[c9][d252][n252];
        end
    endgenerate
    generate 
        localparam integer d253 = 1;
        for (n253 = 0; n253 < 16; n253 = n253 + 1) 
        begin: outbit253
            assign data_11[n253 + d253*16 + c9*28*16] = data_11_array[c9][d253][n253];
        end
    endgenerate
    generate 
        localparam integer d254 = 2;
        for (n254 = 0; n254 < 16; n254 = n254 + 1) 
        begin: outbit254
            assign data_11[n254 + d254*16 + c9*28*16] = data_11_array[c9][d254][n254];
        end
    endgenerate
    generate 
        localparam integer d255 = 3;
        for (n255 = 0; n255 < 16; n255 = n255 + 1) 
        begin: outbit255
            assign data_11[n255 + d255*16 + c9*28*16] = data_11_array[c9][d255][n255];
        end
    endgenerate
    generate 
        localparam integer d256 = 4;
        for (n256 = 0; n256 < 16; n256 = n256 + 1) 
        begin: outbit256
            assign data_11[n256 + d256*16 + c9*28*16] = data_11_array[c9][d256][n256];
        end
    endgenerate
    generate 
        localparam integer d257 = 5;
        for (n257 = 0; n257 < 16; n257 = n257 + 1) 
        begin: outbit257
            assign data_11[n257 + d257*16 + c9*28*16] = data_11_array[c9][d257][n257];
        end
    endgenerate
    generate 
        localparam integer d258 = 6;
        for (n258 = 0; n258 < 16; n258 = n258 + 1) 
        begin: outbit258
            assign data_11[n258 + d258*16 + c9*28*16] = data_11_array[c9][d258][n258];
        end
    endgenerate
    generate 
        localparam integer d259 = 7;
        for (n259 = 0; n259 < 16; n259 = n259 + 1) 
        begin: outbit259
            assign data_11[n259 + d259*16 + c9*28*16] = data_11_array[c9][d259][n259];
        end
    endgenerate
    generate 
        localparam integer d260 = 8;
        for (n260 = 0; n260 < 16; n260 = n260 + 1) 
        begin: outbit260
            assign data_11[n260 + d260*16 + c9*28*16] = data_11_array[c9][d260][n260];
        end
    endgenerate
    generate 
        localparam integer d261 = 9;
        for (n261 = 0; n261 < 16; n261 = n261 + 1) 
        begin: outbit261
            assign data_11[n261 + d261*16 + c9*28*16] = data_11_array[c9][d261][n261];
        end
    endgenerate
    generate 
        localparam integer d262 = 10;
        for (n262 = 0; n262 < 16; n262 = n262 + 1) 
        begin: outbit262
            assign data_11[n262 + d262*16 + c9*28*16] = data_11_array[c9][d262][n262];
        end
    endgenerate
    generate 
        localparam integer d263 = 11;
        for (n263 = 0; n263 < 16; n263 = n263 + 1) 
        begin: outbit263
            assign data_11[n263 + d263*16 + c9*28*16] = data_11_array[c9][d263][n263];
        end
    endgenerate
    generate 
        localparam integer d264 = 12;
        for (n264 = 0; n264 < 16; n264 = n264 + 1) 
        begin: outbit264
            assign data_11[n264 + d264*16 + c9*28*16] = data_11_array[c9][d264][n264];
        end
    endgenerate
    generate 
        localparam integer d265 = 13;
        for (n265 = 0; n265 < 16; n265 = n265 + 1) 
        begin: outbit265
            assign data_11[n265 + d265*16 + c9*28*16] = data_11_array[c9][d265][n265];
        end
    endgenerate
    generate 
        localparam integer d266 = 14;
        for (n266 = 0; n266 < 16; n266 = n266 + 1) 
        begin: outbit266
            assign data_11[n266 + d266*16 + c9*28*16] = data_11_array[c9][d266][n266];
        end
    endgenerate
    generate 
        localparam integer d267 = 15;
        for (n267 = 0; n267 < 16; n267 = n267 + 1) 
        begin: outbit267
            assign data_11[n267 + d267*16 + c9*28*16] = data_11_array[c9][d267][n267];
        end
    endgenerate
    generate 
        localparam integer d268 = 16;
        for (n268 = 0; n268 < 16; n268 = n268 + 1) 
        begin: outbit268
            assign data_11[n268 + d268*16 + c9*28*16] = data_11_array[c9][d268][n268];
        end
    endgenerate
    generate 
        localparam integer d269 = 17;
        for (n269 = 0; n269 < 16; n269 = n269 + 1) 
        begin: outbit269
            assign data_11[n269 + d269*16 + c9*28*16] = data_11_array[c9][d269][n269];
        end
    endgenerate
    generate 
        localparam integer d270 = 18;
        for (n270 = 0; n270 < 16; n270 = n270 + 1) 
        begin: outbit270
            assign data_11[n270 + d270*16 + c9*28*16] = data_11_array[c9][d270][n270];
        end
    endgenerate
    generate 
        localparam integer d271 = 19;
        for (n271 = 0; n271 < 16; n271 = n271 + 1) 
        begin: outbit271
            assign data_11[n271 + d271*16 + c9*28*16] = data_11_array[c9][d271][n271];
        end
    endgenerate
    generate 
        localparam integer d272 = 20;
        for (n272 = 0; n272 < 16; n272 = n272 + 1) 
        begin: outbit272
            assign data_11[n272 + d272*16 + c9*28*16] = data_11_array[c9][d272][n272];
        end
    endgenerate
    generate 
        localparam integer d273 = 21;
        for (n273 = 0; n273 < 16; n273 = n273 + 1) 
        begin: outbit273
            assign data_11[n273 + d273*16 + c9*28*16] = data_11_array[c9][d273][n273];
        end
    endgenerate
    generate 
        localparam integer d274 = 22;
        for (n274 = 0; n274 < 16; n274 = n274 + 1) 
        begin: outbit274
            assign data_11[n274 + d274*16 + c9*28*16] = data_11_array[c9][d274][n274];
        end
    endgenerate
    generate 
        localparam integer d275 = 23;
        for (n275 = 0; n275 < 16; n275 = n275 + 1) 
        begin: outbit275
            assign data_11[n275 + d275*16 + c9*28*16] = data_11_array[c9][d275][n275];
        end
    endgenerate
    generate 
        localparam integer d276 = 24;
        for (n276 = 0; n276 < 16; n276 = n276 + 1) 
        begin: outbit276
            assign data_11[n276 + d276*16 + c9*28*16] = data_11_array[c9][d276][n276];
        end
    endgenerate
    generate 
        localparam integer d277 = 25;
        for (n277 = 0; n277 < 16; n277 = n277 + 1) 
        begin: outbit277
            assign data_11[n277 + d277*16 + c9*28*16] = data_11_array[c9][d277][n277];
        end
    endgenerate
    generate 
        localparam integer d278 = 26;
        for (n278 = 0; n278 < 16; n278 = n278 + 1) 
        begin: outbit278
            assign data_11[n278 + d278*16 + c9*28*16] = data_11_array[c9][d278][n278];
        end
    endgenerate
    generate 
        localparam integer d279 = 27;
        for (n279 = 0; n279 < 16; n279 = n279 + 1) 
        begin: outbit279
            assign data_11[n279 + d279*16 + c9*28*16] = data_11_array[c9][d279][n279];
        end
    endgenerate
    localparam integer c10 = 10;
    generate 
        localparam integer d280 = 0;
        for (n280 = 0; n280 < 16; n280 = n280 + 1) 
        begin: outbit280
            assign data_11[n280 + d280*16 + c10*28*16] = data_11_array[c10][d280][n280];
        end
    endgenerate
    generate 
        localparam integer d281 = 1;
        for (n281 = 0; n281 < 16; n281 = n281 + 1) 
        begin: outbit281
            assign data_11[n281 + d281*16 + c10*28*16] = data_11_array[c10][d281][n281];
        end
    endgenerate
    generate 
        localparam integer d282 = 2;
        for (n282 = 0; n282 < 16; n282 = n282 + 1) 
        begin: outbit282
            assign data_11[n282 + d282*16 + c10*28*16] = data_11_array[c10][d282][n282];
        end
    endgenerate
    generate 
        localparam integer d283 = 3;
        for (n283 = 0; n283 < 16; n283 = n283 + 1) 
        begin: outbit283
            assign data_11[n283 + d283*16 + c10*28*16] = data_11_array[c10][d283][n283];
        end
    endgenerate
    generate 
        localparam integer d284 = 4;
        for (n284 = 0; n284 < 16; n284 = n284 + 1) 
        begin: outbit284
            assign data_11[n284 + d284*16 + c10*28*16] = data_11_array[c10][d284][n284];
        end
    endgenerate
    generate 
        localparam integer d285 = 5;
        for (n285 = 0; n285 < 16; n285 = n285 + 1) 
        begin: outbit285
            assign data_11[n285 + d285*16 + c10*28*16] = data_11_array[c10][d285][n285];
        end
    endgenerate
    generate 
        localparam integer d286 = 6;
        for (n286 = 0; n286 < 16; n286 = n286 + 1) 
        begin: outbit286
            assign data_11[n286 + d286*16 + c10*28*16] = data_11_array[c10][d286][n286];
        end
    endgenerate
    generate 
        localparam integer d287 = 7;
        for (n287 = 0; n287 < 16; n287 = n287 + 1) 
        begin: outbit287
            assign data_11[n287 + d287*16 + c10*28*16] = data_11_array[c10][d287][n287];
        end
    endgenerate
    generate 
        localparam integer d288 = 8;
        for (n288 = 0; n288 < 16; n288 = n288 + 1) 
        begin: outbit288
            assign data_11[n288 + d288*16 + c10*28*16] = data_11_array[c10][d288][n288];
        end
    endgenerate
    generate 
        localparam integer d289 = 9;
        for (n289 = 0; n289 < 16; n289 = n289 + 1) 
        begin: outbit289
            assign data_11[n289 + d289*16 + c10*28*16] = data_11_array[c10][d289][n289];
        end
    endgenerate
    generate 
        localparam integer d290 = 10;
        for (n290 = 0; n290 < 16; n290 = n290 + 1) 
        begin: outbit290
            assign data_11[n290 + d290*16 + c10*28*16] = data_11_array[c10][d290][n290];
        end
    endgenerate
    generate 
        localparam integer d291 = 11;
        for (n291 = 0; n291 < 16; n291 = n291 + 1) 
        begin: outbit291
            assign data_11[n291 + d291*16 + c10*28*16] = data_11_array[c10][d291][n291];
        end
    endgenerate
    generate 
        localparam integer d292 = 12;
        for (n292 = 0; n292 < 16; n292 = n292 + 1) 
        begin: outbit292
            assign data_11[n292 + d292*16 + c10*28*16] = data_11_array[c10][d292][n292];
        end
    endgenerate
    generate 
        localparam integer d293 = 13;
        for (n293 = 0; n293 < 16; n293 = n293 + 1) 
        begin: outbit293
            assign data_11[n293 + d293*16 + c10*28*16] = data_11_array[c10][d293][n293];
        end
    endgenerate
    generate 
        localparam integer d294 = 14;
        for (n294 = 0; n294 < 16; n294 = n294 + 1) 
        begin: outbit294
            assign data_11[n294 + d294*16 + c10*28*16] = data_11_array[c10][d294][n294];
        end
    endgenerate
    generate 
        localparam integer d295 = 15;
        for (n295 = 0; n295 < 16; n295 = n295 + 1) 
        begin: outbit295
            assign data_11[n295 + d295*16 + c10*28*16] = data_11_array[c10][d295][n295];
        end
    endgenerate
    generate 
        localparam integer d296 = 16;
        for (n296 = 0; n296 < 16; n296 = n296 + 1) 
        begin: outbit296
            assign data_11[n296 + d296*16 + c10*28*16] = data_11_array[c10][d296][n296];
        end
    endgenerate
    generate 
        localparam integer d297 = 17;
        for (n297 = 0; n297 < 16; n297 = n297 + 1) 
        begin: outbit297
            assign data_11[n297 + d297*16 + c10*28*16] = data_11_array[c10][d297][n297];
        end
    endgenerate
    generate 
        localparam integer d298 = 18;
        for (n298 = 0; n298 < 16; n298 = n298 + 1) 
        begin: outbit298
            assign data_11[n298 + d298*16 + c10*28*16] = data_11_array[c10][d298][n298];
        end
    endgenerate
    generate 
        localparam integer d299 = 19;
        for (n299 = 0; n299 < 16; n299 = n299 + 1) 
        begin: outbit299
            assign data_11[n299 + d299*16 + c10*28*16] = data_11_array[c10][d299][n299];
        end
    endgenerate
    generate 
        localparam integer d300 = 20;
        for (n300 = 0; n300 < 16; n300 = n300 + 1) 
        begin: outbit300
            assign data_11[n300 + d300*16 + c10*28*16] = data_11_array[c10][d300][n300];
        end
    endgenerate
    generate 
        localparam integer d301 = 21;
        for (n301 = 0; n301 < 16; n301 = n301 + 1) 
        begin: outbit301
            assign data_11[n301 + d301*16 + c10*28*16] = data_11_array[c10][d301][n301];
        end
    endgenerate
    generate 
        localparam integer d302 = 22;
        for (n302 = 0; n302 < 16; n302 = n302 + 1) 
        begin: outbit302
            assign data_11[n302 + d302*16 + c10*28*16] = data_11_array[c10][d302][n302];
        end
    endgenerate
    generate 
        localparam integer d303 = 23;
        for (n303 = 0; n303 < 16; n303 = n303 + 1) 
        begin: outbit303
            assign data_11[n303 + d303*16 + c10*28*16] = data_11_array[c10][d303][n303];
        end
    endgenerate
    generate 
        localparam integer d304 = 24;
        for (n304 = 0; n304 < 16; n304 = n304 + 1) 
        begin: outbit304
            assign data_11[n304 + d304*16 + c10*28*16] = data_11_array[c10][d304][n304];
        end
    endgenerate
    generate 
        localparam integer d305 = 25;
        for (n305 = 0; n305 < 16; n305 = n305 + 1) 
        begin: outbit305
            assign data_11[n305 + d305*16 + c10*28*16] = data_11_array[c10][d305][n305];
        end
    endgenerate
    generate 
        localparam integer d306 = 26;
        for (n306 = 0; n306 < 16; n306 = n306 + 1) 
        begin: outbit306
            assign data_11[n306 + d306*16 + c10*28*16] = data_11_array[c10][d306][n306];
        end
    endgenerate
    generate 
        localparam integer d307 = 27;
        for (n307 = 0; n307 < 16; n307 = n307 + 1) 
        begin: outbit307
            assign data_11[n307 + d307*16 + c10*28*16] = data_11_array[c10][d307][n307];
        end
    endgenerate
    localparam integer c11 = 11;
    generate 
        localparam integer d308 = 0;
        for (n308 = 0; n308 < 16; n308 = n308 + 1) 
        begin: outbit308
            assign data_11[n308 + d308*16 + c11*28*16] = data_11_array[c11][d308][n308];
        end
    endgenerate
    generate 
        localparam integer d309 = 1;
        for (n309 = 0; n309 < 16; n309 = n309 + 1) 
        begin: outbit309
            assign data_11[n309 + d309*16 + c11*28*16] = data_11_array[c11][d309][n309];
        end
    endgenerate
    generate 
        localparam integer d310 = 2;
        for (n310 = 0; n310 < 16; n310 = n310 + 1) 
        begin: outbit310
            assign data_11[n310 + d310*16 + c11*28*16] = data_11_array[c11][d310][n310];
        end
    endgenerate
    generate 
        localparam integer d311 = 3;
        for (n311 = 0; n311 < 16; n311 = n311 + 1) 
        begin: outbit311
            assign data_11[n311 + d311*16 + c11*28*16] = data_11_array[c11][d311][n311];
        end
    endgenerate
    generate 
        localparam integer d312 = 4;
        for (n312 = 0; n312 < 16; n312 = n312 + 1) 
        begin: outbit312
            assign data_11[n312 + d312*16 + c11*28*16] = data_11_array[c11][d312][n312];
        end
    endgenerate
    generate 
        localparam integer d313 = 5;
        for (n313 = 0; n313 < 16; n313 = n313 + 1) 
        begin: outbit313
            assign data_11[n313 + d313*16 + c11*28*16] = data_11_array[c11][d313][n313];
        end
    endgenerate
    generate 
        localparam integer d314 = 6;
        for (n314 = 0; n314 < 16; n314 = n314 + 1) 
        begin: outbit314
            assign data_11[n314 + d314*16 + c11*28*16] = data_11_array[c11][d314][n314];
        end
    endgenerate
    generate 
        localparam integer d315 = 7;
        for (n315 = 0; n315 < 16; n315 = n315 + 1) 
        begin: outbit315
            assign data_11[n315 + d315*16 + c11*28*16] = data_11_array[c11][d315][n315];
        end
    endgenerate
    generate 
        localparam integer d316 = 8;
        for (n316 = 0; n316 < 16; n316 = n316 + 1) 
        begin: outbit316
            assign data_11[n316 + d316*16 + c11*28*16] = data_11_array[c11][d316][n316];
        end
    endgenerate
    generate 
        localparam integer d317 = 9;
        for (n317 = 0; n317 < 16; n317 = n317 + 1) 
        begin: outbit317
            assign data_11[n317 + d317*16 + c11*28*16] = data_11_array[c11][d317][n317];
        end
    endgenerate
    generate 
        localparam integer d318 = 10;
        for (n318 = 0; n318 < 16; n318 = n318 + 1) 
        begin: outbit318
            assign data_11[n318 + d318*16 + c11*28*16] = data_11_array[c11][d318][n318];
        end
    endgenerate
    generate 
        localparam integer d319 = 11;
        for (n319 = 0; n319 < 16; n319 = n319 + 1) 
        begin: outbit319
            assign data_11[n319 + d319*16 + c11*28*16] = data_11_array[c11][d319][n319];
        end
    endgenerate
    generate 
        localparam integer d320 = 12;
        for (n320 = 0; n320 < 16; n320 = n320 + 1) 
        begin: outbit320
            assign data_11[n320 + d320*16 + c11*28*16] = data_11_array[c11][d320][n320];
        end
    endgenerate
    generate 
        localparam integer d321 = 13;
        for (n321 = 0; n321 < 16; n321 = n321 + 1) 
        begin: outbit321
            assign data_11[n321 + d321*16 + c11*28*16] = data_11_array[c11][d321][n321];
        end
    endgenerate
    generate 
        localparam integer d322 = 14;
        for (n322 = 0; n322 < 16; n322 = n322 + 1) 
        begin: outbit322
            assign data_11[n322 + d322*16 + c11*28*16] = data_11_array[c11][d322][n322];
        end
    endgenerate
    generate 
        localparam integer d323 = 15;
        for (n323 = 0; n323 < 16; n323 = n323 + 1) 
        begin: outbit323
            assign data_11[n323 + d323*16 + c11*28*16] = data_11_array[c11][d323][n323];
        end
    endgenerate
    generate 
        localparam integer d324 = 16;
        for (n324 = 0; n324 < 16; n324 = n324 + 1) 
        begin: outbit324
            assign data_11[n324 + d324*16 + c11*28*16] = data_11_array[c11][d324][n324];
        end
    endgenerate
    generate 
        localparam integer d325 = 17;
        for (n325 = 0; n325 < 16; n325 = n325 + 1) 
        begin: outbit325
            assign data_11[n325 + d325*16 + c11*28*16] = data_11_array[c11][d325][n325];
        end
    endgenerate
    generate 
        localparam integer d326 = 18;
        for (n326 = 0; n326 < 16; n326 = n326 + 1) 
        begin: outbit326
            assign data_11[n326 + d326*16 + c11*28*16] = data_11_array[c11][d326][n326];
        end
    endgenerate
    generate 
        localparam integer d327 = 19;
        for (n327 = 0; n327 < 16; n327 = n327 + 1) 
        begin: outbit327
            assign data_11[n327 + d327*16 + c11*28*16] = data_11_array[c11][d327][n327];
        end
    endgenerate
    generate 
        localparam integer d328 = 20;
        for (n328 = 0; n328 < 16; n328 = n328 + 1) 
        begin: outbit328
            assign data_11[n328 + d328*16 + c11*28*16] = data_11_array[c11][d328][n328];
        end
    endgenerate
    generate 
        localparam integer d329 = 21;
        for (n329 = 0; n329 < 16; n329 = n329 + 1) 
        begin: outbit329
            assign data_11[n329 + d329*16 + c11*28*16] = data_11_array[c11][d329][n329];
        end
    endgenerate
    generate 
        localparam integer d330 = 22;
        for (n330 = 0; n330 < 16; n330 = n330 + 1) 
        begin: outbit330
            assign data_11[n330 + d330*16 + c11*28*16] = data_11_array[c11][d330][n330];
        end
    endgenerate
    generate 
        localparam integer d331 = 23;
        for (n331 = 0; n331 < 16; n331 = n331 + 1) 
        begin: outbit331
            assign data_11[n331 + d331*16 + c11*28*16] = data_11_array[c11][d331][n331];
        end
    endgenerate
    generate 
        localparam integer d332 = 24;
        for (n332 = 0; n332 < 16; n332 = n332 + 1) 
        begin: outbit332
            assign data_11[n332 + d332*16 + c11*28*16] = data_11_array[c11][d332][n332];
        end
    endgenerate
    generate 
        localparam integer d333 = 25;
        for (n333 = 0; n333 < 16; n333 = n333 + 1) 
        begin: outbit333
            assign data_11[n333 + d333*16 + c11*28*16] = data_11_array[c11][d333][n333];
        end
    endgenerate
    generate 
        localparam integer d334 = 26;
        for (n334 = 0; n334 < 16; n334 = n334 + 1) 
        begin: outbit334
            assign data_11[n334 + d334*16 + c11*28*16] = data_11_array[c11][d334][n334];
        end
    endgenerate
    generate 
        localparam integer d335 = 27;
        for (n335 = 0; n335 < 16; n335 = n335 + 1) 
        begin: outbit335
            assign data_11[n335 + d335*16 + c11*28*16] = data_11_array[c11][d335][n335];
        end
    endgenerate
    localparam integer c12 = 12;
    generate 
        localparam integer d336 = 0;
        for (n336 = 0; n336 < 16; n336 = n336 + 1) 
        begin: outbit336
            assign data_11[n336 + d336*16 + c12*28*16] = data_11_array[c12][d336][n336];
        end
    endgenerate
    generate 
        localparam integer d337 = 1;
        for (n337 = 0; n337 < 16; n337 = n337 + 1) 
        begin: outbit337
            assign data_11[n337 + d337*16 + c12*28*16] = data_11_array[c12][d337][n337];
        end
    endgenerate
    generate 
        localparam integer d338 = 2;
        for (n338 = 0; n338 < 16; n338 = n338 + 1) 
        begin: outbit338
            assign data_11[n338 + d338*16 + c12*28*16] = data_11_array[c12][d338][n338];
        end
    endgenerate
    generate 
        localparam integer d339 = 3;
        for (n339 = 0; n339 < 16; n339 = n339 + 1) 
        begin: outbit339
            assign data_11[n339 + d339*16 + c12*28*16] = data_11_array[c12][d339][n339];
        end
    endgenerate
    generate 
        localparam integer d340 = 4;
        for (n340 = 0; n340 < 16; n340 = n340 + 1) 
        begin: outbit340
            assign data_11[n340 + d340*16 + c12*28*16] = data_11_array[c12][d340][n340];
        end
    endgenerate
    generate 
        localparam integer d341 = 5;
        for (n341 = 0; n341 < 16; n341 = n341 + 1) 
        begin: outbit341
            assign data_11[n341 + d341*16 + c12*28*16] = data_11_array[c12][d341][n341];
        end
    endgenerate
    generate 
        localparam integer d342 = 6;
        for (n342 = 0; n342 < 16; n342 = n342 + 1) 
        begin: outbit342
            assign data_11[n342 + d342*16 + c12*28*16] = data_11_array[c12][d342][n342];
        end
    endgenerate
    generate 
        localparam integer d343 = 7;
        for (n343 = 0; n343 < 16; n343 = n343 + 1) 
        begin: outbit343
            assign data_11[n343 + d343*16 + c12*28*16] = data_11_array[c12][d343][n343];
        end
    endgenerate
    generate 
        localparam integer d344 = 8;
        for (n344 = 0; n344 < 16; n344 = n344 + 1) 
        begin: outbit344
            assign data_11[n344 + d344*16 + c12*28*16] = data_11_array[c12][d344][n344];
        end
    endgenerate
    generate 
        localparam integer d345 = 9;
        for (n345 = 0; n345 < 16; n345 = n345 + 1) 
        begin: outbit345
            assign data_11[n345 + d345*16 + c12*28*16] = data_11_array[c12][d345][n345];
        end
    endgenerate
    generate 
        localparam integer d346 = 10;
        for (n346 = 0; n346 < 16; n346 = n346 + 1) 
        begin: outbit346
            assign data_11[n346 + d346*16 + c12*28*16] = data_11_array[c12][d346][n346];
        end
    endgenerate
    generate 
        localparam integer d347 = 11;
        for (n347 = 0; n347 < 16; n347 = n347 + 1) 
        begin: outbit347
            assign data_11[n347 + d347*16 + c12*28*16] = data_11_array[c12][d347][n347];
        end
    endgenerate
    generate 
        localparam integer d348 = 12;
        for (n348 = 0; n348 < 16; n348 = n348 + 1) 
        begin: outbit348
            assign data_11[n348 + d348*16 + c12*28*16] = data_11_array[c12][d348][n348];
        end
    endgenerate
    generate 
        localparam integer d349 = 13;
        for (n349 = 0; n349 < 16; n349 = n349 + 1) 
        begin: outbit349
            assign data_11[n349 + d349*16 + c12*28*16] = data_11_array[c12][d349][n349];
        end
    endgenerate
    generate 
        localparam integer d350 = 14;
        for (n350 = 0; n350 < 16; n350 = n350 + 1) 
        begin: outbit350
            assign data_11[n350 + d350*16 + c12*28*16] = data_11_array[c12][d350][n350];
        end
    endgenerate
    generate 
        localparam integer d351 = 15;
        for (n351 = 0; n351 < 16; n351 = n351 + 1) 
        begin: outbit351
            assign data_11[n351 + d351*16 + c12*28*16] = data_11_array[c12][d351][n351];
        end
    endgenerate
    generate 
        localparam integer d352 = 16;
        for (n352 = 0; n352 < 16; n352 = n352 + 1) 
        begin: outbit352
            assign data_11[n352 + d352*16 + c12*28*16] = data_11_array[c12][d352][n352];
        end
    endgenerate
    generate 
        localparam integer d353 = 17;
        for (n353 = 0; n353 < 16; n353 = n353 + 1) 
        begin: outbit353
            assign data_11[n353 + d353*16 + c12*28*16] = data_11_array[c12][d353][n353];
        end
    endgenerate
    generate 
        localparam integer d354 = 18;
        for (n354 = 0; n354 < 16; n354 = n354 + 1) 
        begin: outbit354
            assign data_11[n354 + d354*16 + c12*28*16] = data_11_array[c12][d354][n354];
        end
    endgenerate
    generate 
        localparam integer d355 = 19;
        for (n355 = 0; n355 < 16; n355 = n355 + 1) 
        begin: outbit355
            assign data_11[n355 + d355*16 + c12*28*16] = data_11_array[c12][d355][n355];
        end
    endgenerate
    generate 
        localparam integer d356 = 20;
        for (n356 = 0; n356 < 16; n356 = n356 + 1) 
        begin: outbit356
            assign data_11[n356 + d356*16 + c12*28*16] = data_11_array[c12][d356][n356];
        end
    endgenerate
    generate 
        localparam integer d357 = 21;
        for (n357 = 0; n357 < 16; n357 = n357 + 1) 
        begin: outbit357
            assign data_11[n357 + d357*16 + c12*28*16] = data_11_array[c12][d357][n357];
        end
    endgenerate
    generate 
        localparam integer d358 = 22;
        for (n358 = 0; n358 < 16; n358 = n358 + 1) 
        begin: outbit358
            assign data_11[n358 + d358*16 + c12*28*16] = data_11_array[c12][d358][n358];
        end
    endgenerate
    generate 
        localparam integer d359 = 23;
        for (n359 = 0; n359 < 16; n359 = n359 + 1) 
        begin: outbit359
            assign data_11[n359 + d359*16 + c12*28*16] = data_11_array[c12][d359][n359];
        end
    endgenerate
    generate 
        localparam integer d360 = 24;
        for (n360 = 0; n360 < 16; n360 = n360 + 1) 
        begin: outbit360
            assign data_11[n360 + d360*16 + c12*28*16] = data_11_array[c12][d360][n360];
        end
    endgenerate
    generate 
        localparam integer d361 = 25;
        for (n361 = 0; n361 < 16; n361 = n361 + 1) 
        begin: outbit361
            assign data_11[n361 + d361*16 + c12*28*16] = data_11_array[c12][d361][n361];
        end
    endgenerate
    generate 
        localparam integer d362 = 26;
        for (n362 = 0; n362 < 16; n362 = n362 + 1) 
        begin: outbit362
            assign data_11[n362 + d362*16 + c12*28*16] = data_11_array[c12][d362][n362];
        end
    endgenerate
    generate 
        localparam integer d363 = 27;
        for (n363 = 0; n363 < 16; n363 = n363 + 1) 
        begin: outbit363
            assign data_11[n363 + d363*16 + c12*28*16] = data_11_array[c12][d363][n363];
        end
    endgenerate
    localparam integer c13 = 13;
    generate 
        localparam integer d364 = 0;
        for (n364 = 0; n364 < 16; n364 = n364 + 1) 
        begin: outbit364
            assign data_11[n364 + d364*16 + c13*28*16] = data_11_array[c13][d364][n364];
        end
    endgenerate
    generate 
        localparam integer d365 = 1;
        for (n365 = 0; n365 < 16; n365 = n365 + 1) 
        begin: outbit365
            assign data_11[n365 + d365*16 + c13*28*16] = data_11_array[c13][d365][n365];
        end
    endgenerate
    generate 
        localparam integer d366 = 2;
        for (n366 = 0; n366 < 16; n366 = n366 + 1) 
        begin: outbit366
            assign data_11[n366 + d366*16 + c13*28*16] = data_11_array[c13][d366][n366];
        end
    endgenerate
    generate 
        localparam integer d367 = 3;
        for (n367 = 0; n367 < 16; n367 = n367 + 1) 
        begin: outbit367
            assign data_11[n367 + d367*16 + c13*28*16] = data_11_array[c13][d367][n367];
        end
    endgenerate
    generate 
        localparam integer d368 = 4;
        for (n368 = 0; n368 < 16; n368 = n368 + 1) 
        begin: outbit368
            assign data_11[n368 + d368*16 + c13*28*16] = data_11_array[c13][d368][n368];
        end
    endgenerate
    generate 
        localparam integer d369 = 5;
        for (n369 = 0; n369 < 16; n369 = n369 + 1) 
        begin: outbit369
            assign data_11[n369 + d369*16 + c13*28*16] = data_11_array[c13][d369][n369];
        end
    endgenerate
    generate 
        localparam integer d370 = 6;
        for (n370 = 0; n370 < 16; n370 = n370 + 1) 
        begin: outbit370
            assign data_11[n370 + d370*16 + c13*28*16] = data_11_array[c13][d370][n370];
        end
    endgenerate
    generate 
        localparam integer d371 = 7;
        for (n371 = 0; n371 < 16; n371 = n371 + 1) 
        begin: outbit371
            assign data_11[n371 + d371*16 + c13*28*16] = data_11_array[c13][d371][n371];
        end
    endgenerate
    generate 
        localparam integer d372 = 8;
        for (n372 = 0; n372 < 16; n372 = n372 + 1) 
        begin: outbit372
            assign data_11[n372 + d372*16 + c13*28*16] = data_11_array[c13][d372][n372];
        end
    endgenerate
    generate 
        localparam integer d373 = 9;
        for (n373 = 0; n373 < 16; n373 = n373 + 1) 
        begin: outbit373
            assign data_11[n373 + d373*16 + c13*28*16] = data_11_array[c13][d373][n373];
        end
    endgenerate
    generate 
        localparam integer d374 = 10;
        for (n374 = 0; n374 < 16; n374 = n374 + 1) 
        begin: outbit374
            assign data_11[n374 + d374*16 + c13*28*16] = data_11_array[c13][d374][n374];
        end
    endgenerate
    generate 
        localparam integer d375 = 11;
        for (n375 = 0; n375 < 16; n375 = n375 + 1) 
        begin: outbit375
            assign data_11[n375 + d375*16 + c13*28*16] = data_11_array[c13][d375][n375];
        end
    endgenerate
    generate 
        localparam integer d376 = 12;
        for (n376 = 0; n376 < 16; n376 = n376 + 1) 
        begin: outbit376
            assign data_11[n376 + d376*16 + c13*28*16] = data_11_array[c13][d376][n376];
        end
    endgenerate
    generate 
        localparam integer d377 = 13;
        for (n377 = 0; n377 < 16; n377 = n377 + 1) 
        begin: outbit377
            assign data_11[n377 + d377*16 + c13*28*16] = data_11_array[c13][d377][n377];
        end
    endgenerate
    generate 
        localparam integer d378 = 14;
        for (n378 = 0; n378 < 16; n378 = n378 + 1) 
        begin: outbit378
            assign data_11[n378 + d378*16 + c13*28*16] = data_11_array[c13][d378][n378];
        end
    endgenerate
    generate 
        localparam integer d379 = 15;
        for (n379 = 0; n379 < 16; n379 = n379 + 1) 
        begin: outbit379
            assign data_11[n379 + d379*16 + c13*28*16] = data_11_array[c13][d379][n379];
        end
    endgenerate
    generate 
        localparam integer d380 = 16;
        for (n380 = 0; n380 < 16; n380 = n380 + 1) 
        begin: outbit380
            assign data_11[n380 + d380*16 + c13*28*16] = data_11_array[c13][d380][n380];
        end
    endgenerate
    generate 
        localparam integer d381 = 17;
        for (n381 = 0; n381 < 16; n381 = n381 + 1) 
        begin: outbit381
            assign data_11[n381 + d381*16 + c13*28*16] = data_11_array[c13][d381][n381];
        end
    endgenerate
    generate 
        localparam integer d382 = 18;
        for (n382 = 0; n382 < 16; n382 = n382 + 1) 
        begin: outbit382
            assign data_11[n382 + d382*16 + c13*28*16] = data_11_array[c13][d382][n382];
        end
    endgenerate
    generate 
        localparam integer d383 = 19;
        for (n383 = 0; n383 < 16; n383 = n383 + 1) 
        begin: outbit383
            assign data_11[n383 + d383*16 + c13*28*16] = data_11_array[c13][d383][n383];
        end
    endgenerate
    generate 
        localparam integer d384 = 20;
        for (n384 = 0; n384 < 16; n384 = n384 + 1) 
        begin: outbit384
            assign data_11[n384 + d384*16 + c13*28*16] = data_11_array[c13][d384][n384];
        end
    endgenerate
    generate 
        localparam integer d385 = 21;
        for (n385 = 0; n385 < 16; n385 = n385 + 1) 
        begin: outbit385
            assign data_11[n385 + d385*16 + c13*28*16] = data_11_array[c13][d385][n385];
        end
    endgenerate
    generate 
        localparam integer d386 = 22;
        for (n386 = 0; n386 < 16; n386 = n386 + 1) 
        begin: outbit386
            assign data_11[n386 + d386*16 + c13*28*16] = data_11_array[c13][d386][n386];
        end
    endgenerate
    generate 
        localparam integer d387 = 23;
        for (n387 = 0; n387 < 16; n387 = n387 + 1) 
        begin: outbit387
            assign data_11[n387 + d387*16 + c13*28*16] = data_11_array[c13][d387][n387];
        end
    endgenerate
    generate 
        localparam integer d388 = 24;
        for (n388 = 0; n388 < 16; n388 = n388 + 1) 
        begin: outbit388
            assign data_11[n388 + d388*16 + c13*28*16] = data_11_array[c13][d388][n388];
        end
    endgenerate
    generate 
        localparam integer d389 = 25;
        for (n389 = 0; n389 < 16; n389 = n389 + 1) 
        begin: outbit389
            assign data_11[n389 + d389*16 + c13*28*16] = data_11_array[c13][d389][n389];
        end
    endgenerate
    generate 
        localparam integer d390 = 26;
        for (n390 = 0; n390 < 16; n390 = n390 + 1) 
        begin: outbit390
            assign data_11[n390 + d390*16 + c13*28*16] = data_11_array[c13][d390][n390];
        end
    endgenerate
    generate 
        localparam integer d391 = 27;
        for (n391 = 0; n391 < 16; n391 = n391 + 1) 
        begin: outbit391
            assign data_11[n391 + d391*16 + c13*28*16] = data_11_array[c13][d391][n391];
        end
    endgenerate
    localparam integer c14 = 14;
    generate 
        localparam integer d392 = 0;
        for (n392 = 0; n392 < 16; n392 = n392 + 1) 
        begin: outbit392
            assign data_11[n392 + d392*16 + c14*28*16] = data_11_array[c14][d392][n392];
        end
    endgenerate
    generate 
        localparam integer d393 = 1;
        for (n393 = 0; n393 < 16; n393 = n393 + 1) 
        begin: outbit393
            assign data_11[n393 + d393*16 + c14*28*16] = data_11_array[c14][d393][n393];
        end
    endgenerate
    generate 
        localparam integer d394 = 2;
        for (n394 = 0; n394 < 16; n394 = n394 + 1) 
        begin: outbit394
            assign data_11[n394 + d394*16 + c14*28*16] = data_11_array[c14][d394][n394];
        end
    endgenerate
    generate 
        localparam integer d395 = 3;
        for (n395 = 0; n395 < 16; n395 = n395 + 1) 
        begin: outbit395
            assign data_11[n395 + d395*16 + c14*28*16] = data_11_array[c14][d395][n395];
        end
    endgenerate
    generate 
        localparam integer d396 = 4;
        for (n396 = 0; n396 < 16; n396 = n396 + 1) 
        begin: outbit396
            assign data_11[n396 + d396*16 + c14*28*16] = data_11_array[c14][d396][n396];
        end
    endgenerate
    generate 
        localparam integer d397 = 5;
        for (n397 = 0; n397 < 16; n397 = n397 + 1) 
        begin: outbit397
            assign data_11[n397 + d397*16 + c14*28*16] = data_11_array[c14][d397][n397];
        end
    endgenerate
    generate 
        localparam integer d398 = 6;
        for (n398 = 0; n398 < 16; n398 = n398 + 1) 
        begin: outbit398
            assign data_11[n398 + d398*16 + c14*28*16] = data_11_array[c14][d398][n398];
        end
    endgenerate
    generate 
        localparam integer d399 = 7;
        for (n399 = 0; n399 < 16; n399 = n399 + 1) 
        begin: outbit399
            assign data_11[n399 + d399*16 + c14*28*16] = data_11_array[c14][d399][n399];
        end
    endgenerate
    generate 
        localparam integer d400 = 8;
        for (n400 = 0; n400 < 16; n400 = n400 + 1) 
        begin: outbit400
            assign data_11[n400 + d400*16 + c14*28*16] = data_11_array[c14][d400][n400];
        end
    endgenerate
    generate 
        localparam integer d401 = 9;
        for (n401 = 0; n401 < 16; n401 = n401 + 1) 
        begin: outbit401
            assign data_11[n401 + d401*16 + c14*28*16] = data_11_array[c14][d401][n401];
        end
    endgenerate
    generate 
        localparam integer d402 = 10;
        for (n402 = 0; n402 < 16; n402 = n402 + 1) 
        begin: outbit402
            assign data_11[n402 + d402*16 + c14*28*16] = data_11_array[c14][d402][n402];
        end
    endgenerate
    generate 
        localparam integer d403 = 11;
        for (n403 = 0; n403 < 16; n403 = n403 + 1) 
        begin: outbit403
            assign data_11[n403 + d403*16 + c14*28*16] = data_11_array[c14][d403][n403];
        end
    endgenerate
    generate 
        localparam integer d404 = 12;
        for (n404 = 0; n404 < 16; n404 = n404 + 1) 
        begin: outbit404
            assign data_11[n404 + d404*16 + c14*28*16] = data_11_array[c14][d404][n404];
        end
    endgenerate
    generate 
        localparam integer d405 = 13;
        for (n405 = 0; n405 < 16; n405 = n405 + 1) 
        begin: outbit405
            assign data_11[n405 + d405*16 + c14*28*16] = data_11_array[c14][d405][n405];
        end
    endgenerate
    generate 
        localparam integer d406 = 14;
        for (n406 = 0; n406 < 16; n406 = n406 + 1) 
        begin: outbit406
            assign data_11[n406 + d406*16 + c14*28*16] = data_11_array[c14][d406][n406];
        end
    endgenerate
    generate 
        localparam integer d407 = 15;
        for (n407 = 0; n407 < 16; n407 = n407 + 1) 
        begin: outbit407
            assign data_11[n407 + d407*16 + c14*28*16] = data_11_array[c14][d407][n407];
        end
    endgenerate
    generate 
        localparam integer d408 = 16;
        for (n408 = 0; n408 < 16; n408 = n408 + 1) 
        begin: outbit408
            assign data_11[n408 + d408*16 + c14*28*16] = data_11_array[c14][d408][n408];
        end
    endgenerate
    generate 
        localparam integer d409 = 17;
        for (n409 = 0; n409 < 16; n409 = n409 + 1) 
        begin: outbit409
            assign data_11[n409 + d409*16 + c14*28*16] = data_11_array[c14][d409][n409];
        end
    endgenerate
    generate 
        localparam integer d410 = 18;
        for (n410 = 0; n410 < 16; n410 = n410 + 1) 
        begin: outbit410
            assign data_11[n410 + d410*16 + c14*28*16] = data_11_array[c14][d410][n410];
        end
    endgenerate
    generate 
        localparam integer d411 = 19;
        for (n411 = 0; n411 < 16; n411 = n411 + 1) 
        begin: outbit411
            assign data_11[n411 + d411*16 + c14*28*16] = data_11_array[c14][d411][n411];
        end
    endgenerate
    generate 
        localparam integer d412 = 20;
        for (n412 = 0; n412 < 16; n412 = n412 + 1) 
        begin: outbit412
            assign data_11[n412 + d412*16 + c14*28*16] = data_11_array[c14][d412][n412];
        end
    endgenerate
    generate 
        localparam integer d413 = 21;
        for (n413 = 0; n413 < 16; n413 = n413 + 1) 
        begin: outbit413
            assign data_11[n413 + d413*16 + c14*28*16] = data_11_array[c14][d413][n413];
        end
    endgenerate
    generate 
        localparam integer d414 = 22;
        for (n414 = 0; n414 < 16; n414 = n414 + 1) 
        begin: outbit414
            assign data_11[n414 + d414*16 + c14*28*16] = data_11_array[c14][d414][n414];
        end
    endgenerate
    generate 
        localparam integer d415 = 23;
        for (n415 = 0; n415 < 16; n415 = n415 + 1) 
        begin: outbit415
            assign data_11[n415 + d415*16 + c14*28*16] = data_11_array[c14][d415][n415];
        end
    endgenerate
    generate 
        localparam integer d416 = 24;
        for (n416 = 0; n416 < 16; n416 = n416 + 1) 
        begin: outbit416
            assign data_11[n416 + d416*16 + c14*28*16] = data_11_array[c14][d416][n416];
        end
    endgenerate
    generate 
        localparam integer d417 = 25;
        for (n417 = 0; n417 < 16; n417 = n417 + 1) 
        begin: outbit417
            assign data_11[n417 + d417*16 + c14*28*16] = data_11_array[c14][d417][n417];
        end
    endgenerate
    generate 
        localparam integer d418 = 26;
        for (n418 = 0; n418 < 16; n418 = n418 + 1) 
        begin: outbit418
            assign data_11[n418 + d418*16 + c14*28*16] = data_11_array[c14][d418][n418];
        end
    endgenerate
    generate 
        localparam integer d419 = 27;
        for (n419 = 0; n419 < 16; n419 = n419 + 1) 
        begin: outbit419
            assign data_11[n419 + d419*16 + c14*28*16] = data_11_array[c14][d419][n419];
        end
    endgenerate
    localparam integer c15 = 15;
    generate 
        localparam integer d420 = 0;
        for (n420 = 0; n420 < 16; n420 = n420 + 1) 
        begin: outbit420
            assign data_11[n420 + d420*16 + c15*28*16] = data_11_array[c15][d420][n420];
        end
    endgenerate
    generate 
        localparam integer d421 = 1;
        for (n421 = 0; n421 < 16; n421 = n421 + 1) 
        begin: outbit421
            assign data_11[n421 + d421*16 + c15*28*16] = data_11_array[c15][d421][n421];
        end
    endgenerate
    generate 
        localparam integer d422 = 2;
        for (n422 = 0; n422 < 16; n422 = n422 + 1) 
        begin: outbit422
            assign data_11[n422 + d422*16 + c15*28*16] = data_11_array[c15][d422][n422];
        end
    endgenerate
    generate 
        localparam integer d423 = 3;
        for (n423 = 0; n423 < 16; n423 = n423 + 1) 
        begin: outbit423
            assign data_11[n423 + d423*16 + c15*28*16] = data_11_array[c15][d423][n423];
        end
    endgenerate
    generate 
        localparam integer d424 = 4;
        for (n424 = 0; n424 < 16; n424 = n424 + 1) 
        begin: outbit424
            assign data_11[n424 + d424*16 + c15*28*16] = data_11_array[c15][d424][n424];
        end
    endgenerate
    generate 
        localparam integer d425 = 5;
        for (n425 = 0; n425 < 16; n425 = n425 + 1) 
        begin: outbit425
            assign data_11[n425 + d425*16 + c15*28*16] = data_11_array[c15][d425][n425];
        end
    endgenerate
    generate 
        localparam integer d426 = 6;
        for (n426 = 0; n426 < 16; n426 = n426 + 1) 
        begin: outbit426
            assign data_11[n426 + d426*16 + c15*28*16] = data_11_array[c15][d426][n426];
        end
    endgenerate
    generate 
        localparam integer d427 = 7;
        for (n427 = 0; n427 < 16; n427 = n427 + 1) 
        begin: outbit427
            assign data_11[n427 + d427*16 + c15*28*16] = data_11_array[c15][d427][n427];
        end
    endgenerate
    generate 
        localparam integer d428 = 8;
        for (n428 = 0; n428 < 16; n428 = n428 + 1) 
        begin: outbit428
            assign data_11[n428 + d428*16 + c15*28*16] = data_11_array[c15][d428][n428];
        end
    endgenerate
    generate 
        localparam integer d429 = 9;
        for (n429 = 0; n429 < 16; n429 = n429 + 1) 
        begin: outbit429
            assign data_11[n429 + d429*16 + c15*28*16] = data_11_array[c15][d429][n429];
        end
    endgenerate
    generate 
        localparam integer d430 = 10;
        for (n430 = 0; n430 < 16; n430 = n430 + 1) 
        begin: outbit430
            assign data_11[n430 + d430*16 + c15*28*16] = data_11_array[c15][d430][n430];
        end
    endgenerate
    generate 
        localparam integer d431 = 11;
        for (n431 = 0; n431 < 16; n431 = n431 + 1) 
        begin: outbit431
            assign data_11[n431 + d431*16 + c15*28*16] = data_11_array[c15][d431][n431];
        end
    endgenerate
    generate 
        localparam integer d432 = 12;
        for (n432 = 0; n432 < 16; n432 = n432 + 1) 
        begin: outbit432
            assign data_11[n432 + d432*16 + c15*28*16] = data_11_array[c15][d432][n432];
        end
    endgenerate
    generate 
        localparam integer d433 = 13;
        for (n433 = 0; n433 < 16; n433 = n433 + 1) 
        begin: outbit433
            assign data_11[n433 + d433*16 + c15*28*16] = data_11_array[c15][d433][n433];
        end
    endgenerate
    generate 
        localparam integer d434 = 14;
        for (n434 = 0; n434 < 16; n434 = n434 + 1) 
        begin: outbit434
            assign data_11[n434 + d434*16 + c15*28*16] = data_11_array[c15][d434][n434];
        end
    endgenerate
    generate 
        localparam integer d435 = 15;
        for (n435 = 0; n435 < 16; n435 = n435 + 1) 
        begin: outbit435
            assign data_11[n435 + d435*16 + c15*28*16] = data_11_array[c15][d435][n435];
        end
    endgenerate
    generate 
        localparam integer d436 = 16;
        for (n436 = 0; n436 < 16; n436 = n436 + 1) 
        begin: outbit436
            assign data_11[n436 + d436*16 + c15*28*16] = data_11_array[c15][d436][n436];
        end
    endgenerate
    generate 
        localparam integer d437 = 17;
        for (n437 = 0; n437 < 16; n437 = n437 + 1) 
        begin: outbit437
            assign data_11[n437 + d437*16 + c15*28*16] = data_11_array[c15][d437][n437];
        end
    endgenerate
    generate 
        localparam integer d438 = 18;
        for (n438 = 0; n438 < 16; n438 = n438 + 1) 
        begin: outbit438
            assign data_11[n438 + d438*16 + c15*28*16] = data_11_array[c15][d438][n438];
        end
    endgenerate
    generate 
        localparam integer d439 = 19;
        for (n439 = 0; n439 < 16; n439 = n439 + 1) 
        begin: outbit439
            assign data_11[n439 + d439*16 + c15*28*16] = data_11_array[c15][d439][n439];
        end
    endgenerate
    generate 
        localparam integer d440 = 20;
        for (n440 = 0; n440 < 16; n440 = n440 + 1) 
        begin: outbit440
            assign data_11[n440 + d440*16 + c15*28*16] = data_11_array[c15][d440][n440];
        end
    endgenerate
    generate 
        localparam integer d441 = 21;
        for (n441 = 0; n441 < 16; n441 = n441 + 1) 
        begin: outbit441
            assign data_11[n441 + d441*16 + c15*28*16] = data_11_array[c15][d441][n441];
        end
    endgenerate
    generate 
        localparam integer d442 = 22;
        for (n442 = 0; n442 < 16; n442 = n442 + 1) 
        begin: outbit442
            assign data_11[n442 + d442*16 + c15*28*16] = data_11_array[c15][d442][n442];
        end
    endgenerate
    generate 
        localparam integer d443 = 23;
        for (n443 = 0; n443 < 16; n443 = n443 + 1) 
        begin: outbit443
            assign data_11[n443 + d443*16 + c15*28*16] = data_11_array[c15][d443][n443];
        end
    endgenerate
    generate 
        localparam integer d444 = 24;
        for (n444 = 0; n444 < 16; n444 = n444 + 1) 
        begin: outbit444
            assign data_11[n444 + d444*16 + c15*28*16] = data_11_array[c15][d444][n444];
        end
    endgenerate
    generate 
        localparam integer d445 = 25;
        for (n445 = 0; n445 < 16; n445 = n445 + 1) 
        begin: outbit445
            assign data_11[n445 + d445*16 + c15*28*16] = data_11_array[c15][d445][n445];
        end
    endgenerate
    generate 
        localparam integer d446 = 26;
        for (n446 = 0; n446 < 16; n446 = n446 + 1) 
        begin: outbit446
            assign data_11[n446 + d446*16 + c15*28*16] = data_11_array[c15][d446][n446];
        end
    endgenerate
    generate 
        localparam integer d447 = 27;
        for (n447 = 0; n447 < 16; n447 = n447 + 1) 
        begin: outbit447
            assign data_11[n447 + d447*16 + c15*28*16] = data_11_array[c15][d447][n447];
        end
    endgenerate
    localparam integer c16 = 16;
    generate 
        localparam integer d448 = 0;
        for (n448 = 0; n448 < 16; n448 = n448 + 1) 
        begin: outbit448
            assign data_11[n448 + d448*16 + c16*28*16] = data_11_array[c16][d448][n448];
        end
    endgenerate
    generate 
        localparam integer d449 = 1;
        for (n449 = 0; n449 < 16; n449 = n449 + 1) 
        begin: outbit449
            assign data_11[n449 + d449*16 + c16*28*16] = data_11_array[c16][d449][n449];
        end
    endgenerate
    generate 
        localparam integer d450 = 2;
        for (n450 = 0; n450 < 16; n450 = n450 + 1) 
        begin: outbit450
            assign data_11[n450 + d450*16 + c16*28*16] = data_11_array[c16][d450][n450];
        end
    endgenerate
    generate 
        localparam integer d451 = 3;
        for (n451 = 0; n451 < 16; n451 = n451 + 1) 
        begin: outbit451
            assign data_11[n451 + d451*16 + c16*28*16] = data_11_array[c16][d451][n451];
        end
    endgenerate
    generate 
        localparam integer d452 = 4;
        for (n452 = 0; n452 < 16; n452 = n452 + 1) 
        begin: outbit452
            assign data_11[n452 + d452*16 + c16*28*16] = data_11_array[c16][d452][n452];
        end
    endgenerate
    generate 
        localparam integer d453 = 5;
        for (n453 = 0; n453 < 16; n453 = n453 + 1) 
        begin: outbit453
            assign data_11[n453 + d453*16 + c16*28*16] = data_11_array[c16][d453][n453];
        end
    endgenerate
    generate 
        localparam integer d454 = 6;
        for (n454 = 0; n454 < 16; n454 = n454 + 1) 
        begin: outbit454
            assign data_11[n454 + d454*16 + c16*28*16] = data_11_array[c16][d454][n454];
        end
    endgenerate
    generate 
        localparam integer d455 = 7;
        for (n455 = 0; n455 < 16; n455 = n455 + 1) 
        begin: outbit455
            assign data_11[n455 + d455*16 + c16*28*16] = data_11_array[c16][d455][n455];
        end
    endgenerate
    generate 
        localparam integer d456 = 8;
        for (n456 = 0; n456 < 16; n456 = n456 + 1) 
        begin: outbit456
            assign data_11[n456 + d456*16 + c16*28*16] = data_11_array[c16][d456][n456];
        end
    endgenerate
    generate 
        localparam integer d457 = 9;
        for (n457 = 0; n457 < 16; n457 = n457 + 1) 
        begin: outbit457
            assign data_11[n457 + d457*16 + c16*28*16] = data_11_array[c16][d457][n457];
        end
    endgenerate
    generate 
        localparam integer d458 = 10;
        for (n458 = 0; n458 < 16; n458 = n458 + 1) 
        begin: outbit458
            assign data_11[n458 + d458*16 + c16*28*16] = data_11_array[c16][d458][n458];
        end
    endgenerate
    generate 
        localparam integer d459 = 11;
        for (n459 = 0; n459 < 16; n459 = n459 + 1) 
        begin: outbit459
            assign data_11[n459 + d459*16 + c16*28*16] = data_11_array[c16][d459][n459];
        end
    endgenerate
    generate 
        localparam integer d460 = 12;
        for (n460 = 0; n460 < 16; n460 = n460 + 1) 
        begin: outbit460
            assign data_11[n460 + d460*16 + c16*28*16] = data_11_array[c16][d460][n460];
        end
    endgenerate
    generate 
        localparam integer d461 = 13;
        for (n461 = 0; n461 < 16; n461 = n461 + 1) 
        begin: outbit461
            assign data_11[n461 + d461*16 + c16*28*16] = data_11_array[c16][d461][n461];
        end
    endgenerate
    generate 
        localparam integer d462 = 14;
        for (n462 = 0; n462 < 16; n462 = n462 + 1) 
        begin: outbit462
            assign data_11[n462 + d462*16 + c16*28*16] = data_11_array[c16][d462][n462];
        end
    endgenerate
    generate 
        localparam integer d463 = 15;
        for (n463 = 0; n463 < 16; n463 = n463 + 1) 
        begin: outbit463
            assign data_11[n463 + d463*16 + c16*28*16] = data_11_array[c16][d463][n463];
        end
    endgenerate
    generate 
        localparam integer d464 = 16;
        for (n464 = 0; n464 < 16; n464 = n464 + 1) 
        begin: outbit464
            assign data_11[n464 + d464*16 + c16*28*16] = data_11_array[c16][d464][n464];
        end
    endgenerate
    generate 
        localparam integer d465 = 17;
        for (n465 = 0; n465 < 16; n465 = n465 + 1) 
        begin: outbit465
            assign data_11[n465 + d465*16 + c16*28*16] = data_11_array[c16][d465][n465];
        end
    endgenerate
    generate 
        localparam integer d466 = 18;
        for (n466 = 0; n466 < 16; n466 = n466 + 1) 
        begin: outbit466
            assign data_11[n466 + d466*16 + c16*28*16] = data_11_array[c16][d466][n466];
        end
    endgenerate
    generate 
        localparam integer d467 = 19;
        for (n467 = 0; n467 < 16; n467 = n467 + 1) 
        begin: outbit467
            assign data_11[n467 + d467*16 + c16*28*16] = data_11_array[c16][d467][n467];
        end
    endgenerate
    generate 
        localparam integer d468 = 20;
        for (n468 = 0; n468 < 16; n468 = n468 + 1) 
        begin: outbit468
            assign data_11[n468 + d468*16 + c16*28*16] = data_11_array[c16][d468][n468];
        end
    endgenerate
    generate 
        localparam integer d469 = 21;
        for (n469 = 0; n469 < 16; n469 = n469 + 1) 
        begin: outbit469
            assign data_11[n469 + d469*16 + c16*28*16] = data_11_array[c16][d469][n469];
        end
    endgenerate
    generate 
        localparam integer d470 = 22;
        for (n470 = 0; n470 < 16; n470 = n470 + 1) 
        begin: outbit470
            assign data_11[n470 + d470*16 + c16*28*16] = data_11_array[c16][d470][n470];
        end
    endgenerate
    generate 
        localparam integer d471 = 23;
        for (n471 = 0; n471 < 16; n471 = n471 + 1) 
        begin: outbit471
            assign data_11[n471 + d471*16 + c16*28*16] = data_11_array[c16][d471][n471];
        end
    endgenerate
    generate 
        localparam integer d472 = 24;
        for (n472 = 0; n472 < 16; n472 = n472 + 1) 
        begin: outbit472
            assign data_11[n472 + d472*16 + c16*28*16] = data_11_array[c16][d472][n472];
        end
    endgenerate
    generate 
        localparam integer d473 = 25;
        for (n473 = 0; n473 < 16; n473 = n473 + 1) 
        begin: outbit473
            assign data_11[n473 + d473*16 + c16*28*16] = data_11_array[c16][d473][n473];
        end
    endgenerate
    generate 
        localparam integer d474 = 26;
        for (n474 = 0; n474 < 16; n474 = n474 + 1) 
        begin: outbit474
            assign data_11[n474 + d474*16 + c16*28*16] = data_11_array[c16][d474][n474];
        end
    endgenerate
    generate 
        localparam integer d475 = 27;
        for (n475 = 0; n475 < 16; n475 = n475 + 1) 
        begin: outbit475
            assign data_11[n475 + d475*16 + c16*28*16] = data_11_array[c16][d475][n475];
        end
    endgenerate
    localparam integer c17 = 17;
    generate 
        localparam integer d476 = 0;
        for (n476 = 0; n476 < 16; n476 = n476 + 1) 
        begin: outbit476
            assign data_11[n476 + d476*16 + c17*28*16] = data_11_array[c17][d476][n476];
        end
    endgenerate
    generate 
        localparam integer d477 = 1;
        for (n477 = 0; n477 < 16; n477 = n477 + 1) 
        begin: outbit477
            assign data_11[n477 + d477*16 + c17*28*16] = data_11_array[c17][d477][n477];
        end
    endgenerate
    generate 
        localparam integer d478 = 2;
        for (n478 = 0; n478 < 16; n478 = n478 + 1) 
        begin: outbit478
            assign data_11[n478 + d478*16 + c17*28*16] = data_11_array[c17][d478][n478];
        end
    endgenerate
    generate 
        localparam integer d479 = 3;
        for (n479 = 0; n479 < 16; n479 = n479 + 1) 
        begin: outbit479
            assign data_11[n479 + d479*16 + c17*28*16] = data_11_array[c17][d479][n479];
        end
    endgenerate
    generate 
        localparam integer d480 = 4;
        for (n480 = 0; n480 < 16; n480 = n480 + 1) 
        begin: outbit480
            assign data_11[n480 + d480*16 + c17*28*16] = data_11_array[c17][d480][n480];
        end
    endgenerate
    generate 
        localparam integer d481 = 5;
        for (n481 = 0; n481 < 16; n481 = n481 + 1) 
        begin: outbit481
            assign data_11[n481 + d481*16 + c17*28*16] = data_11_array[c17][d481][n481];
        end
    endgenerate
    generate 
        localparam integer d482 = 6;
        for (n482 = 0; n482 < 16; n482 = n482 + 1) 
        begin: outbit482
            assign data_11[n482 + d482*16 + c17*28*16] = data_11_array[c17][d482][n482];
        end
    endgenerate
    generate 
        localparam integer d483 = 7;
        for (n483 = 0; n483 < 16; n483 = n483 + 1) 
        begin: outbit483
            assign data_11[n483 + d483*16 + c17*28*16] = data_11_array[c17][d483][n483];
        end
    endgenerate
    generate 
        localparam integer d484 = 8;
        for (n484 = 0; n484 < 16; n484 = n484 + 1) 
        begin: outbit484
            assign data_11[n484 + d484*16 + c17*28*16] = data_11_array[c17][d484][n484];
        end
    endgenerate
    generate 
        localparam integer d485 = 9;
        for (n485 = 0; n485 < 16; n485 = n485 + 1) 
        begin: outbit485
            assign data_11[n485 + d485*16 + c17*28*16] = data_11_array[c17][d485][n485];
        end
    endgenerate
    generate 
        localparam integer d486 = 10;
        for (n486 = 0; n486 < 16; n486 = n486 + 1) 
        begin: outbit486
            assign data_11[n486 + d486*16 + c17*28*16] = data_11_array[c17][d486][n486];
        end
    endgenerate
    generate 
        localparam integer d487 = 11;
        for (n487 = 0; n487 < 16; n487 = n487 + 1) 
        begin: outbit487
            assign data_11[n487 + d487*16 + c17*28*16] = data_11_array[c17][d487][n487];
        end
    endgenerate
    generate 
        localparam integer d488 = 12;
        for (n488 = 0; n488 < 16; n488 = n488 + 1) 
        begin: outbit488
            assign data_11[n488 + d488*16 + c17*28*16] = data_11_array[c17][d488][n488];
        end
    endgenerate
    generate 
        localparam integer d489 = 13;
        for (n489 = 0; n489 < 16; n489 = n489 + 1) 
        begin: outbit489
            assign data_11[n489 + d489*16 + c17*28*16] = data_11_array[c17][d489][n489];
        end
    endgenerate
    generate 
        localparam integer d490 = 14;
        for (n490 = 0; n490 < 16; n490 = n490 + 1) 
        begin: outbit490
            assign data_11[n490 + d490*16 + c17*28*16] = data_11_array[c17][d490][n490];
        end
    endgenerate
    generate 
        localparam integer d491 = 15;
        for (n491 = 0; n491 < 16; n491 = n491 + 1) 
        begin: outbit491
            assign data_11[n491 + d491*16 + c17*28*16] = data_11_array[c17][d491][n491];
        end
    endgenerate
    generate 
        localparam integer d492 = 16;
        for (n492 = 0; n492 < 16; n492 = n492 + 1) 
        begin: outbit492
            assign data_11[n492 + d492*16 + c17*28*16] = data_11_array[c17][d492][n492];
        end
    endgenerate
    generate 
        localparam integer d493 = 17;
        for (n493 = 0; n493 < 16; n493 = n493 + 1) 
        begin: outbit493
            assign data_11[n493 + d493*16 + c17*28*16] = data_11_array[c17][d493][n493];
        end
    endgenerate
    generate 
        localparam integer d494 = 18;
        for (n494 = 0; n494 < 16; n494 = n494 + 1) 
        begin: outbit494
            assign data_11[n494 + d494*16 + c17*28*16] = data_11_array[c17][d494][n494];
        end
    endgenerate
    generate 
        localparam integer d495 = 19;
        for (n495 = 0; n495 < 16; n495 = n495 + 1) 
        begin: outbit495
            assign data_11[n495 + d495*16 + c17*28*16] = data_11_array[c17][d495][n495];
        end
    endgenerate
    generate 
        localparam integer d496 = 20;
        for (n496 = 0; n496 < 16; n496 = n496 + 1) 
        begin: outbit496
            assign data_11[n496 + d496*16 + c17*28*16] = data_11_array[c17][d496][n496];
        end
    endgenerate
    generate 
        localparam integer d497 = 21;
        for (n497 = 0; n497 < 16; n497 = n497 + 1) 
        begin: outbit497
            assign data_11[n497 + d497*16 + c17*28*16] = data_11_array[c17][d497][n497];
        end
    endgenerate
    generate 
        localparam integer d498 = 22;
        for (n498 = 0; n498 < 16; n498 = n498 + 1) 
        begin: outbit498
            assign data_11[n498 + d498*16 + c17*28*16] = data_11_array[c17][d498][n498];
        end
    endgenerate
    generate 
        localparam integer d499 = 23;
        for (n499 = 0; n499 < 16; n499 = n499 + 1) 
        begin: outbit499
            assign data_11[n499 + d499*16 + c17*28*16] = data_11_array[c17][d499][n499];
        end
    endgenerate
    generate 
        localparam integer d500 = 24;
        for (n500 = 0; n500 < 16; n500 = n500 + 1) 
        begin: outbit500
            assign data_11[n500 + d500*16 + c17*28*16] = data_11_array[c17][d500][n500];
        end
    endgenerate
    generate 
        localparam integer d501 = 25;
        for (n501 = 0; n501 < 16; n501 = n501 + 1) 
        begin: outbit501
            assign data_11[n501 + d501*16 + c17*28*16] = data_11_array[c17][d501][n501];
        end
    endgenerate
    generate 
        localparam integer d502 = 26;
        for (n502 = 0; n502 < 16; n502 = n502 + 1) 
        begin: outbit502
            assign data_11[n502 + d502*16 + c17*28*16] = data_11_array[c17][d502][n502];
        end
    endgenerate
    generate 
        localparam integer d503 = 27;
        for (n503 = 0; n503 < 16; n503 = n503 + 1) 
        begin: outbit503
            assign data_11[n503 + d503*16 + c17*28*16] = data_11_array[c17][d503][n503];
        end
    endgenerate
    localparam integer c18 = 18;
    generate 
        localparam integer d504 = 0;
        for (n504 = 0; n504 < 16; n504 = n504 + 1) 
        begin: outbit504
            assign data_11[n504 + d504*16 + c18*28*16] = data_11_array[c18][d504][n504];
        end
    endgenerate
    generate 
        localparam integer d505 = 1;
        for (n505 = 0; n505 < 16; n505 = n505 + 1) 
        begin: outbit505
            assign data_11[n505 + d505*16 + c18*28*16] = data_11_array[c18][d505][n505];
        end
    endgenerate
    generate 
        localparam integer d506 = 2;
        for (n506 = 0; n506 < 16; n506 = n506 + 1) 
        begin: outbit506
            assign data_11[n506 + d506*16 + c18*28*16] = data_11_array[c18][d506][n506];
        end
    endgenerate
    generate 
        localparam integer d507 = 3;
        for (n507 = 0; n507 < 16; n507 = n507 + 1) 
        begin: outbit507
            assign data_11[n507 + d507*16 + c18*28*16] = data_11_array[c18][d507][n507];
        end
    endgenerate
    generate 
        localparam integer d508 = 4;
        for (n508 = 0; n508 < 16; n508 = n508 + 1) 
        begin: outbit508
            assign data_11[n508 + d508*16 + c18*28*16] = data_11_array[c18][d508][n508];
        end
    endgenerate
    generate 
        localparam integer d509 = 5;
        for (n509 = 0; n509 < 16; n509 = n509 + 1) 
        begin: outbit509
            assign data_11[n509 + d509*16 + c18*28*16] = data_11_array[c18][d509][n509];
        end
    endgenerate
    generate 
        localparam integer d510 = 6;
        for (n510 = 0; n510 < 16; n510 = n510 + 1) 
        begin: outbit510
            assign data_11[n510 + d510*16 + c18*28*16] = data_11_array[c18][d510][n510];
        end
    endgenerate
    generate 
        localparam integer d511 = 7;
        for (n511 = 0; n511 < 16; n511 = n511 + 1) 
        begin: outbit511
            assign data_11[n511 + d511*16 + c18*28*16] = data_11_array[c18][d511][n511];
        end
    endgenerate
    generate 
        localparam integer d512 = 8;
        for (n512 = 0; n512 < 16; n512 = n512 + 1) 
        begin: outbit512
            assign data_11[n512 + d512*16 + c18*28*16] = data_11_array[c18][d512][n512];
        end
    endgenerate
    generate 
        localparam integer d513 = 9;
        for (n513 = 0; n513 < 16; n513 = n513 + 1) 
        begin: outbit513
            assign data_11[n513 + d513*16 + c18*28*16] = data_11_array[c18][d513][n513];
        end
    endgenerate
    generate 
        localparam integer d514 = 10;
        for (n514 = 0; n514 < 16; n514 = n514 + 1) 
        begin: outbit514
            assign data_11[n514 + d514*16 + c18*28*16] = data_11_array[c18][d514][n514];
        end
    endgenerate
    generate 
        localparam integer d515 = 11;
        for (n515 = 0; n515 < 16; n515 = n515 + 1) 
        begin: outbit515
            assign data_11[n515 + d515*16 + c18*28*16] = data_11_array[c18][d515][n515];
        end
    endgenerate
    generate 
        localparam integer d516 = 12;
        for (n516 = 0; n516 < 16; n516 = n516 + 1) 
        begin: outbit516
            assign data_11[n516 + d516*16 + c18*28*16] = data_11_array[c18][d516][n516];
        end
    endgenerate
    generate 
        localparam integer d517 = 13;
        for (n517 = 0; n517 < 16; n517 = n517 + 1) 
        begin: outbit517
            assign data_11[n517 + d517*16 + c18*28*16] = data_11_array[c18][d517][n517];
        end
    endgenerate
    generate 
        localparam integer d518 = 14;
        for (n518 = 0; n518 < 16; n518 = n518 + 1) 
        begin: outbit518
            assign data_11[n518 + d518*16 + c18*28*16] = data_11_array[c18][d518][n518];
        end
    endgenerate
    generate 
        localparam integer d519 = 15;
        for (n519 = 0; n519 < 16; n519 = n519 + 1) 
        begin: outbit519
            assign data_11[n519 + d519*16 + c18*28*16] = data_11_array[c18][d519][n519];
        end
    endgenerate
    generate 
        localparam integer d520 = 16;
        for (n520 = 0; n520 < 16; n520 = n520 + 1) 
        begin: outbit520
            assign data_11[n520 + d520*16 + c18*28*16] = data_11_array[c18][d520][n520];
        end
    endgenerate
    generate 
        localparam integer d521 = 17;
        for (n521 = 0; n521 < 16; n521 = n521 + 1) 
        begin: outbit521
            assign data_11[n521 + d521*16 + c18*28*16] = data_11_array[c18][d521][n521];
        end
    endgenerate
    generate 
        localparam integer d522 = 18;
        for (n522 = 0; n522 < 16; n522 = n522 + 1) 
        begin: outbit522
            assign data_11[n522 + d522*16 + c18*28*16] = data_11_array[c18][d522][n522];
        end
    endgenerate
    generate 
        localparam integer d523 = 19;
        for (n523 = 0; n523 < 16; n523 = n523 + 1) 
        begin: outbit523
            assign data_11[n523 + d523*16 + c18*28*16] = data_11_array[c18][d523][n523];
        end
    endgenerate
    generate 
        localparam integer d524 = 20;
        for (n524 = 0; n524 < 16; n524 = n524 + 1) 
        begin: outbit524
            assign data_11[n524 + d524*16 + c18*28*16] = data_11_array[c18][d524][n524];
        end
    endgenerate
    generate 
        localparam integer d525 = 21;
        for (n525 = 0; n525 < 16; n525 = n525 + 1) 
        begin: outbit525
            assign data_11[n525 + d525*16 + c18*28*16] = data_11_array[c18][d525][n525];
        end
    endgenerate
    generate 
        localparam integer d526 = 22;
        for (n526 = 0; n526 < 16; n526 = n526 + 1) 
        begin: outbit526
            assign data_11[n526 + d526*16 + c18*28*16] = data_11_array[c18][d526][n526];
        end
    endgenerate
    generate 
        localparam integer d527 = 23;
        for (n527 = 0; n527 < 16; n527 = n527 + 1) 
        begin: outbit527
            assign data_11[n527 + d527*16 + c18*28*16] = data_11_array[c18][d527][n527];
        end
    endgenerate
    generate 
        localparam integer d528 = 24;
        for (n528 = 0; n528 < 16; n528 = n528 + 1) 
        begin: outbit528
            assign data_11[n528 + d528*16 + c18*28*16] = data_11_array[c18][d528][n528];
        end
    endgenerate
    generate 
        localparam integer d529 = 25;
        for (n529 = 0; n529 < 16; n529 = n529 + 1) 
        begin: outbit529
            assign data_11[n529 + d529*16 + c18*28*16] = data_11_array[c18][d529][n529];
        end
    endgenerate
    generate 
        localparam integer d530 = 26;
        for (n530 = 0; n530 < 16; n530 = n530 + 1) 
        begin: outbit530
            assign data_11[n530 + d530*16 + c18*28*16] = data_11_array[c18][d530][n530];
        end
    endgenerate
    generate 
        localparam integer d531 = 27;
        for (n531 = 0; n531 < 16; n531 = n531 + 1) 
        begin: outbit531
            assign data_11[n531 + d531*16 + c18*28*16] = data_11_array[c18][d531][n531];
        end
    endgenerate
    localparam integer c19 = 19;
    generate 
        localparam integer d532 = 0;
        for (n532 = 0; n532 < 16; n532 = n532 + 1) 
        begin: outbit532
            assign data_11[n532 + d532*16 + c19*28*16] = data_11_array[c19][d532][n532];
        end
    endgenerate
    generate 
        localparam integer d533 = 1;
        for (n533 = 0; n533 < 16; n533 = n533 + 1) 
        begin: outbit533
            assign data_11[n533 + d533*16 + c19*28*16] = data_11_array[c19][d533][n533];
        end
    endgenerate
    generate 
        localparam integer d534 = 2;
        for (n534 = 0; n534 < 16; n534 = n534 + 1) 
        begin: outbit534
            assign data_11[n534 + d534*16 + c19*28*16] = data_11_array[c19][d534][n534];
        end
    endgenerate
    generate 
        localparam integer d535 = 3;
        for (n535 = 0; n535 < 16; n535 = n535 + 1) 
        begin: outbit535
            assign data_11[n535 + d535*16 + c19*28*16] = data_11_array[c19][d535][n535];
        end
    endgenerate
    generate 
        localparam integer d536 = 4;
        for (n536 = 0; n536 < 16; n536 = n536 + 1) 
        begin: outbit536
            assign data_11[n536 + d536*16 + c19*28*16] = data_11_array[c19][d536][n536];
        end
    endgenerate
    generate 
        localparam integer d537 = 5;
        for (n537 = 0; n537 < 16; n537 = n537 + 1) 
        begin: outbit537
            assign data_11[n537 + d537*16 + c19*28*16] = data_11_array[c19][d537][n537];
        end
    endgenerate
    generate 
        localparam integer d538 = 6;
        for (n538 = 0; n538 < 16; n538 = n538 + 1) 
        begin: outbit538
            assign data_11[n538 + d538*16 + c19*28*16] = data_11_array[c19][d538][n538];
        end
    endgenerate
    generate 
        localparam integer d539 = 7;
        for (n539 = 0; n539 < 16; n539 = n539 + 1) 
        begin: outbit539
            assign data_11[n539 + d539*16 + c19*28*16] = data_11_array[c19][d539][n539];
        end
    endgenerate
    generate 
        localparam integer d540 = 8;
        for (n540 = 0; n540 < 16; n540 = n540 + 1) 
        begin: outbit540
            assign data_11[n540 + d540*16 + c19*28*16] = data_11_array[c19][d540][n540];
        end
    endgenerate
    generate 
        localparam integer d541 = 9;
        for (n541 = 0; n541 < 16; n541 = n541 + 1) 
        begin: outbit541
            assign data_11[n541 + d541*16 + c19*28*16] = data_11_array[c19][d541][n541];
        end
    endgenerate
    generate 
        localparam integer d542 = 10;
        for (n542 = 0; n542 < 16; n542 = n542 + 1) 
        begin: outbit542
            assign data_11[n542 + d542*16 + c19*28*16] = data_11_array[c19][d542][n542];
        end
    endgenerate
    generate 
        localparam integer d543 = 11;
        for (n543 = 0; n543 < 16; n543 = n543 + 1) 
        begin: outbit543
            assign data_11[n543 + d543*16 + c19*28*16] = data_11_array[c19][d543][n543];
        end
    endgenerate
    generate 
        localparam integer d544 = 12;
        for (n544 = 0; n544 < 16; n544 = n544 + 1) 
        begin: outbit544
            assign data_11[n544 + d544*16 + c19*28*16] = data_11_array[c19][d544][n544];
        end
    endgenerate
    generate 
        localparam integer d545 = 13;
        for (n545 = 0; n545 < 16; n545 = n545 + 1) 
        begin: outbit545
            assign data_11[n545 + d545*16 + c19*28*16] = data_11_array[c19][d545][n545];
        end
    endgenerate
    generate 
        localparam integer d546 = 14;
        for (n546 = 0; n546 < 16; n546 = n546 + 1) 
        begin: outbit546
            assign data_11[n546 + d546*16 + c19*28*16] = data_11_array[c19][d546][n546];
        end
    endgenerate
    generate 
        localparam integer d547 = 15;
        for (n547 = 0; n547 < 16; n547 = n547 + 1) 
        begin: outbit547
            assign data_11[n547 + d547*16 + c19*28*16] = data_11_array[c19][d547][n547];
        end
    endgenerate
    generate 
        localparam integer d548 = 16;
        for (n548 = 0; n548 < 16; n548 = n548 + 1) 
        begin: outbit548
            assign data_11[n548 + d548*16 + c19*28*16] = data_11_array[c19][d548][n548];
        end
    endgenerate
    generate 
        localparam integer d549 = 17;
        for (n549 = 0; n549 < 16; n549 = n549 + 1) 
        begin: outbit549
            assign data_11[n549 + d549*16 + c19*28*16] = data_11_array[c19][d549][n549];
        end
    endgenerate
    generate 
        localparam integer d550 = 18;
        for (n550 = 0; n550 < 16; n550 = n550 + 1) 
        begin: outbit550
            assign data_11[n550 + d550*16 + c19*28*16] = data_11_array[c19][d550][n550];
        end
    endgenerate
    generate 
        localparam integer d551 = 19;
        for (n551 = 0; n551 < 16; n551 = n551 + 1) 
        begin: outbit551
            assign data_11[n551 + d551*16 + c19*28*16] = data_11_array[c19][d551][n551];
        end
    endgenerate
    generate 
        localparam integer d552 = 20;
        for (n552 = 0; n552 < 16; n552 = n552 + 1) 
        begin: outbit552
            assign data_11[n552 + d552*16 + c19*28*16] = data_11_array[c19][d552][n552];
        end
    endgenerate
    generate 
        localparam integer d553 = 21;
        for (n553 = 0; n553 < 16; n553 = n553 + 1) 
        begin: outbit553
            assign data_11[n553 + d553*16 + c19*28*16] = data_11_array[c19][d553][n553];
        end
    endgenerate
    generate 
        localparam integer d554 = 22;
        for (n554 = 0; n554 < 16; n554 = n554 + 1) 
        begin: outbit554
            assign data_11[n554 + d554*16 + c19*28*16] = data_11_array[c19][d554][n554];
        end
    endgenerate
    generate 
        localparam integer d555 = 23;
        for (n555 = 0; n555 < 16; n555 = n555 + 1) 
        begin: outbit555
            assign data_11[n555 + d555*16 + c19*28*16] = data_11_array[c19][d555][n555];
        end
    endgenerate
    generate 
        localparam integer d556 = 24;
        for (n556 = 0; n556 < 16; n556 = n556 + 1) 
        begin: outbit556
            assign data_11[n556 + d556*16 + c19*28*16] = data_11_array[c19][d556][n556];
        end
    endgenerate
    generate 
        localparam integer d557 = 25;
        for (n557 = 0; n557 < 16; n557 = n557 + 1) 
        begin: outbit557
            assign data_11[n557 + d557*16 + c19*28*16] = data_11_array[c19][d557][n557];
        end
    endgenerate
    generate 
        localparam integer d558 = 26;
        for (n558 = 0; n558 < 16; n558 = n558 + 1) 
        begin: outbit558
            assign data_11[n558 + d558*16 + c19*28*16] = data_11_array[c19][d558][n558];
        end
    endgenerate
    generate 
        localparam integer d559 = 27;
        for (n559 = 0; n559 < 16; n559 = n559 + 1) 
        begin: outbit559
            assign data_11[n559 + d559*16 + c19*28*16] = data_11_array[c19][d559][n559];
        end
    endgenerate
    localparam integer c20 = 20;
    generate 
        localparam integer d560 = 0;
        for (n560 = 0; n560 < 16; n560 = n560 + 1) 
        begin: outbit560
            assign data_11[n560 + d560*16 + c20*28*16] = data_11_array[c20][d560][n560];
        end
    endgenerate
    generate 
        localparam integer d561 = 1;
        for (n561 = 0; n561 < 16; n561 = n561 + 1) 
        begin: outbit561
            assign data_11[n561 + d561*16 + c20*28*16] = data_11_array[c20][d561][n561];
        end
    endgenerate
    generate 
        localparam integer d562 = 2;
        for (n562 = 0; n562 < 16; n562 = n562 + 1) 
        begin: outbit562
            assign data_11[n562 + d562*16 + c20*28*16] = data_11_array[c20][d562][n562];
        end
    endgenerate
    generate 
        localparam integer d563 = 3;
        for (n563 = 0; n563 < 16; n563 = n563 + 1) 
        begin: outbit563
            assign data_11[n563 + d563*16 + c20*28*16] = data_11_array[c20][d563][n563];
        end
    endgenerate
    generate 
        localparam integer d564 = 4;
        for (n564 = 0; n564 < 16; n564 = n564 + 1) 
        begin: outbit564
            assign data_11[n564 + d564*16 + c20*28*16] = data_11_array[c20][d564][n564];
        end
    endgenerate
    generate 
        localparam integer d565 = 5;
        for (n565 = 0; n565 < 16; n565 = n565 + 1) 
        begin: outbit565
            assign data_11[n565 + d565*16 + c20*28*16] = data_11_array[c20][d565][n565];
        end
    endgenerate
    generate 
        localparam integer d566 = 6;
        for (n566 = 0; n566 < 16; n566 = n566 + 1) 
        begin: outbit566
            assign data_11[n566 + d566*16 + c20*28*16] = data_11_array[c20][d566][n566];
        end
    endgenerate
    generate 
        localparam integer d567 = 7;
        for (n567 = 0; n567 < 16; n567 = n567 + 1) 
        begin: outbit567
            assign data_11[n567 + d567*16 + c20*28*16] = data_11_array[c20][d567][n567];
        end
    endgenerate
    generate 
        localparam integer d568 = 8;
        for (n568 = 0; n568 < 16; n568 = n568 + 1) 
        begin: outbit568
            assign data_11[n568 + d568*16 + c20*28*16] = data_11_array[c20][d568][n568];
        end
    endgenerate
    generate 
        localparam integer d569 = 9;
        for (n569 = 0; n569 < 16; n569 = n569 + 1) 
        begin: outbit569
            assign data_11[n569 + d569*16 + c20*28*16] = data_11_array[c20][d569][n569];
        end
    endgenerate
    generate 
        localparam integer d570 = 10;
        for (n570 = 0; n570 < 16; n570 = n570 + 1) 
        begin: outbit570
            assign data_11[n570 + d570*16 + c20*28*16] = data_11_array[c20][d570][n570];
        end
    endgenerate
    generate 
        localparam integer d571 = 11;
        for (n571 = 0; n571 < 16; n571 = n571 + 1) 
        begin: outbit571
            assign data_11[n571 + d571*16 + c20*28*16] = data_11_array[c20][d571][n571];
        end
    endgenerate
    generate 
        localparam integer d572 = 12;
        for (n572 = 0; n572 < 16; n572 = n572 + 1) 
        begin: outbit572
            assign data_11[n572 + d572*16 + c20*28*16] = data_11_array[c20][d572][n572];
        end
    endgenerate
    generate 
        localparam integer d573 = 13;
        for (n573 = 0; n573 < 16; n573 = n573 + 1) 
        begin: outbit573
            assign data_11[n573 + d573*16 + c20*28*16] = data_11_array[c20][d573][n573];
        end
    endgenerate
    generate 
        localparam integer d574 = 14;
        for (n574 = 0; n574 < 16; n574 = n574 + 1) 
        begin: outbit574
            assign data_11[n574 + d574*16 + c20*28*16] = data_11_array[c20][d574][n574];
        end
    endgenerate
    generate 
        localparam integer d575 = 15;
        for (n575 = 0; n575 < 16; n575 = n575 + 1) 
        begin: outbit575
            assign data_11[n575 + d575*16 + c20*28*16] = data_11_array[c20][d575][n575];
        end
    endgenerate
    generate 
        localparam integer d576 = 16;
        for (n576 = 0; n576 < 16; n576 = n576 + 1) 
        begin: outbit576
            assign data_11[n576 + d576*16 + c20*28*16] = data_11_array[c20][d576][n576];
        end
    endgenerate
    generate 
        localparam integer d577 = 17;
        for (n577 = 0; n577 < 16; n577 = n577 + 1) 
        begin: outbit577
            assign data_11[n577 + d577*16 + c20*28*16] = data_11_array[c20][d577][n577];
        end
    endgenerate
    generate 
        localparam integer d578 = 18;
        for (n578 = 0; n578 < 16; n578 = n578 + 1) 
        begin: outbit578
            assign data_11[n578 + d578*16 + c20*28*16] = data_11_array[c20][d578][n578];
        end
    endgenerate
    generate 
        localparam integer d579 = 19;
        for (n579 = 0; n579 < 16; n579 = n579 + 1) 
        begin: outbit579
            assign data_11[n579 + d579*16 + c20*28*16] = data_11_array[c20][d579][n579];
        end
    endgenerate
    generate 
        localparam integer d580 = 20;
        for (n580 = 0; n580 < 16; n580 = n580 + 1) 
        begin: outbit580
            assign data_11[n580 + d580*16 + c20*28*16] = data_11_array[c20][d580][n580];
        end
    endgenerate
    generate 
        localparam integer d581 = 21;
        for (n581 = 0; n581 < 16; n581 = n581 + 1) 
        begin: outbit581
            assign data_11[n581 + d581*16 + c20*28*16] = data_11_array[c20][d581][n581];
        end
    endgenerate
    generate 
        localparam integer d582 = 22;
        for (n582 = 0; n582 < 16; n582 = n582 + 1) 
        begin: outbit582
            assign data_11[n582 + d582*16 + c20*28*16] = data_11_array[c20][d582][n582];
        end
    endgenerate
    generate 
        localparam integer d583 = 23;
        for (n583 = 0; n583 < 16; n583 = n583 + 1) 
        begin: outbit583
            assign data_11[n583 + d583*16 + c20*28*16] = data_11_array[c20][d583][n583];
        end
    endgenerate
    generate 
        localparam integer d584 = 24;
        for (n584 = 0; n584 < 16; n584 = n584 + 1) 
        begin: outbit584
            assign data_11[n584 + d584*16 + c20*28*16] = data_11_array[c20][d584][n584];
        end
    endgenerate
    generate 
        localparam integer d585 = 25;
        for (n585 = 0; n585 < 16; n585 = n585 + 1) 
        begin: outbit585
            assign data_11[n585 + d585*16 + c20*28*16] = data_11_array[c20][d585][n585];
        end
    endgenerate
    generate 
        localparam integer d586 = 26;
        for (n586 = 0; n586 < 16; n586 = n586 + 1) 
        begin: outbit586
            assign data_11[n586 + d586*16 + c20*28*16] = data_11_array[c20][d586][n586];
        end
    endgenerate
    generate 
        localparam integer d587 = 27;
        for (n587 = 0; n587 < 16; n587 = n587 + 1) 
        begin: outbit587
            assign data_11[n587 + d587*16 + c20*28*16] = data_11_array[c20][d587][n587];
        end
    endgenerate
    localparam integer c21 = 21;
    generate 
        localparam integer d588 = 0;
        for (n588 = 0; n588 < 16; n588 = n588 + 1) 
        begin: outbit588
            assign data_11[n588 + d588*16 + c21*28*16] = data_11_array[c21][d588][n588];
        end
    endgenerate
    generate 
        localparam integer d589 = 1;
        for (n589 = 0; n589 < 16; n589 = n589 + 1) 
        begin: outbit589
            assign data_11[n589 + d589*16 + c21*28*16] = data_11_array[c21][d589][n589];
        end
    endgenerate
    generate 
        localparam integer d590 = 2;
        for (n590 = 0; n590 < 16; n590 = n590 + 1) 
        begin: outbit590
            assign data_11[n590 + d590*16 + c21*28*16] = data_11_array[c21][d590][n590];
        end
    endgenerate
    generate 
        localparam integer d591 = 3;
        for (n591 = 0; n591 < 16; n591 = n591 + 1) 
        begin: outbit591
            assign data_11[n591 + d591*16 + c21*28*16] = data_11_array[c21][d591][n591];
        end
    endgenerate
    generate 
        localparam integer d592 = 4;
        for (n592 = 0; n592 < 16; n592 = n592 + 1) 
        begin: outbit592
            assign data_11[n592 + d592*16 + c21*28*16] = data_11_array[c21][d592][n592];
        end
    endgenerate
    generate 
        localparam integer d593 = 5;
        for (n593 = 0; n593 < 16; n593 = n593 + 1) 
        begin: outbit593
            assign data_11[n593 + d593*16 + c21*28*16] = data_11_array[c21][d593][n593];
        end
    endgenerate
    generate 
        localparam integer d594 = 6;
        for (n594 = 0; n594 < 16; n594 = n594 + 1) 
        begin: outbit594
            assign data_11[n594 + d594*16 + c21*28*16] = data_11_array[c21][d594][n594];
        end
    endgenerate
    generate 
        localparam integer d595 = 7;
        for (n595 = 0; n595 < 16; n595 = n595 + 1) 
        begin: outbit595
            assign data_11[n595 + d595*16 + c21*28*16] = data_11_array[c21][d595][n595];
        end
    endgenerate
    generate 
        localparam integer d596 = 8;
        for (n596 = 0; n596 < 16; n596 = n596 + 1) 
        begin: outbit596
            assign data_11[n596 + d596*16 + c21*28*16] = data_11_array[c21][d596][n596];
        end
    endgenerate
    generate 
        localparam integer d597 = 9;
        for (n597 = 0; n597 < 16; n597 = n597 + 1) 
        begin: outbit597
            assign data_11[n597 + d597*16 + c21*28*16] = data_11_array[c21][d597][n597];
        end
    endgenerate
    generate 
        localparam integer d598 = 10;
        for (n598 = 0; n598 < 16; n598 = n598 + 1) 
        begin: outbit598
            assign data_11[n598 + d598*16 + c21*28*16] = data_11_array[c21][d598][n598];
        end
    endgenerate
    generate 
        localparam integer d599 = 11;
        for (n599 = 0; n599 < 16; n599 = n599 + 1) 
        begin: outbit599
            assign data_11[n599 + d599*16 + c21*28*16] = data_11_array[c21][d599][n599];
        end
    endgenerate
    generate 
        localparam integer d600 = 12;
        for (n600 = 0; n600 < 16; n600 = n600 + 1) 
        begin: outbit600
            assign data_11[n600 + d600*16 + c21*28*16] = data_11_array[c21][d600][n600];
        end
    endgenerate
    generate 
        localparam integer d601 = 13;
        for (n601 = 0; n601 < 16; n601 = n601 + 1) 
        begin: outbit601
            assign data_11[n601 + d601*16 + c21*28*16] = data_11_array[c21][d601][n601];
        end
    endgenerate
    generate 
        localparam integer d602 = 14;
        for (n602 = 0; n602 < 16; n602 = n602 + 1) 
        begin: outbit602
            assign data_11[n602 + d602*16 + c21*28*16] = data_11_array[c21][d602][n602];
        end
    endgenerate
    generate 
        localparam integer d603 = 15;
        for (n603 = 0; n603 < 16; n603 = n603 + 1) 
        begin: outbit603
            assign data_11[n603 + d603*16 + c21*28*16] = data_11_array[c21][d603][n603];
        end
    endgenerate
    generate 
        localparam integer d604 = 16;
        for (n604 = 0; n604 < 16; n604 = n604 + 1) 
        begin: outbit604
            assign data_11[n604 + d604*16 + c21*28*16] = data_11_array[c21][d604][n604];
        end
    endgenerate
    generate 
        localparam integer d605 = 17;
        for (n605 = 0; n605 < 16; n605 = n605 + 1) 
        begin: outbit605
            assign data_11[n605 + d605*16 + c21*28*16] = data_11_array[c21][d605][n605];
        end
    endgenerate
    generate 
        localparam integer d606 = 18;
        for (n606 = 0; n606 < 16; n606 = n606 + 1) 
        begin: outbit606
            assign data_11[n606 + d606*16 + c21*28*16] = data_11_array[c21][d606][n606];
        end
    endgenerate
    generate 
        localparam integer d607 = 19;
        for (n607 = 0; n607 < 16; n607 = n607 + 1) 
        begin: outbit607
            assign data_11[n607 + d607*16 + c21*28*16] = data_11_array[c21][d607][n607];
        end
    endgenerate
    generate 
        localparam integer d608 = 20;
        for (n608 = 0; n608 < 16; n608 = n608 + 1) 
        begin: outbit608
            assign data_11[n608 + d608*16 + c21*28*16] = data_11_array[c21][d608][n608];
        end
    endgenerate
    generate 
        localparam integer d609 = 21;
        for (n609 = 0; n609 < 16; n609 = n609 + 1) 
        begin: outbit609
            assign data_11[n609 + d609*16 + c21*28*16] = data_11_array[c21][d609][n609];
        end
    endgenerate
    generate 
        localparam integer d610 = 22;
        for (n610 = 0; n610 < 16; n610 = n610 + 1) 
        begin: outbit610
            assign data_11[n610 + d610*16 + c21*28*16] = data_11_array[c21][d610][n610];
        end
    endgenerate
    generate 
        localparam integer d611 = 23;
        for (n611 = 0; n611 < 16; n611 = n611 + 1) 
        begin: outbit611
            assign data_11[n611 + d611*16 + c21*28*16] = data_11_array[c21][d611][n611];
        end
    endgenerate
    generate 
        localparam integer d612 = 24;
        for (n612 = 0; n612 < 16; n612 = n612 + 1) 
        begin: outbit612
            assign data_11[n612 + d612*16 + c21*28*16] = data_11_array[c21][d612][n612];
        end
    endgenerate
    generate 
        localparam integer d613 = 25;
        for (n613 = 0; n613 < 16; n613 = n613 + 1) 
        begin: outbit613
            assign data_11[n613 + d613*16 + c21*28*16] = data_11_array[c21][d613][n613];
        end
    endgenerate
    generate 
        localparam integer d614 = 26;
        for (n614 = 0; n614 < 16; n614 = n614 + 1) 
        begin: outbit614
            assign data_11[n614 + d614*16 + c21*28*16] = data_11_array[c21][d614][n614];
        end
    endgenerate
    generate 
        localparam integer d615 = 27;
        for (n615 = 0; n615 < 16; n615 = n615 + 1) 
        begin: outbit615
            assign data_11[n615 + d615*16 + c21*28*16] = data_11_array[c21][d615][n615];
        end
    endgenerate
    localparam integer c22 = 22;
    generate 
        localparam integer d616 = 0;
        for (n616 = 0; n616 < 16; n616 = n616 + 1) 
        begin: outbit616
            assign data_11[n616 + d616*16 + c22*28*16] = data_11_array[c22][d616][n616];
        end
    endgenerate
    generate 
        localparam integer d617 = 1;
        for (n617 = 0; n617 < 16; n617 = n617 + 1) 
        begin: outbit617
            assign data_11[n617 + d617*16 + c22*28*16] = data_11_array[c22][d617][n617];
        end
    endgenerate
    generate 
        localparam integer d618 = 2;
        for (n618 = 0; n618 < 16; n618 = n618 + 1) 
        begin: outbit618
            assign data_11[n618 + d618*16 + c22*28*16] = data_11_array[c22][d618][n618];
        end
    endgenerate
    generate 
        localparam integer d619 = 3;
        for (n619 = 0; n619 < 16; n619 = n619 + 1) 
        begin: outbit619
            assign data_11[n619 + d619*16 + c22*28*16] = data_11_array[c22][d619][n619];
        end
    endgenerate
    generate 
        localparam integer d620 = 4;
        for (n620 = 0; n620 < 16; n620 = n620 + 1) 
        begin: outbit620
            assign data_11[n620 + d620*16 + c22*28*16] = data_11_array[c22][d620][n620];
        end
    endgenerate
    generate 
        localparam integer d621 = 5;
        for (n621 = 0; n621 < 16; n621 = n621 + 1) 
        begin: outbit621
            assign data_11[n621 + d621*16 + c22*28*16] = data_11_array[c22][d621][n621];
        end
    endgenerate
    generate 
        localparam integer d622 = 6;
        for (n622 = 0; n622 < 16; n622 = n622 + 1) 
        begin: outbit622
            assign data_11[n622 + d622*16 + c22*28*16] = data_11_array[c22][d622][n622];
        end
    endgenerate
    generate 
        localparam integer d623 = 7;
        for (n623 = 0; n623 < 16; n623 = n623 + 1) 
        begin: outbit623
            assign data_11[n623 + d623*16 + c22*28*16] = data_11_array[c22][d623][n623];
        end
    endgenerate
    generate 
        localparam integer d624 = 8;
        for (n624 = 0; n624 < 16; n624 = n624 + 1) 
        begin: outbit624
            assign data_11[n624 + d624*16 + c22*28*16] = data_11_array[c22][d624][n624];
        end
    endgenerate
    generate 
        localparam integer d625 = 9;
        for (n625 = 0; n625 < 16; n625 = n625 + 1) 
        begin: outbit625
            assign data_11[n625 + d625*16 + c22*28*16] = data_11_array[c22][d625][n625];
        end
    endgenerate
    generate 
        localparam integer d626 = 10;
        for (n626 = 0; n626 < 16; n626 = n626 + 1) 
        begin: outbit626
            assign data_11[n626 + d626*16 + c22*28*16] = data_11_array[c22][d626][n626];
        end
    endgenerate
    generate 
        localparam integer d627 = 11;
        for (n627 = 0; n627 < 16; n627 = n627 + 1) 
        begin: outbit627
            assign data_11[n627 + d627*16 + c22*28*16] = data_11_array[c22][d627][n627];
        end
    endgenerate
    generate 
        localparam integer d628 = 12;
        for (n628 = 0; n628 < 16; n628 = n628 + 1) 
        begin: outbit628
            assign data_11[n628 + d628*16 + c22*28*16] = data_11_array[c22][d628][n628];
        end
    endgenerate
    generate 
        localparam integer d629 = 13;
        for (n629 = 0; n629 < 16; n629 = n629 + 1) 
        begin: outbit629
            assign data_11[n629 + d629*16 + c22*28*16] = data_11_array[c22][d629][n629];
        end
    endgenerate
    generate 
        localparam integer d630 = 14;
        for (n630 = 0; n630 < 16; n630 = n630 + 1) 
        begin: outbit630
            assign data_11[n630 + d630*16 + c22*28*16] = data_11_array[c22][d630][n630];
        end
    endgenerate
    generate 
        localparam integer d631 = 15;
        for (n631 = 0; n631 < 16; n631 = n631 + 1) 
        begin: outbit631
            assign data_11[n631 + d631*16 + c22*28*16] = data_11_array[c22][d631][n631];
        end
    endgenerate
    generate 
        localparam integer d632 = 16;
        for (n632 = 0; n632 < 16; n632 = n632 + 1) 
        begin: outbit632
            assign data_11[n632 + d632*16 + c22*28*16] = data_11_array[c22][d632][n632];
        end
    endgenerate
    generate 
        localparam integer d633 = 17;
        for (n633 = 0; n633 < 16; n633 = n633 + 1) 
        begin: outbit633
            assign data_11[n633 + d633*16 + c22*28*16] = data_11_array[c22][d633][n633];
        end
    endgenerate
    generate 
        localparam integer d634 = 18;
        for (n634 = 0; n634 < 16; n634 = n634 + 1) 
        begin: outbit634
            assign data_11[n634 + d634*16 + c22*28*16] = data_11_array[c22][d634][n634];
        end
    endgenerate
    generate 
        localparam integer d635 = 19;
        for (n635 = 0; n635 < 16; n635 = n635 + 1) 
        begin: outbit635
            assign data_11[n635 + d635*16 + c22*28*16] = data_11_array[c22][d635][n635];
        end
    endgenerate
    generate 
        localparam integer d636 = 20;
        for (n636 = 0; n636 < 16; n636 = n636 + 1) 
        begin: outbit636
            assign data_11[n636 + d636*16 + c22*28*16] = data_11_array[c22][d636][n636];
        end
    endgenerate
    generate 
        localparam integer d637 = 21;
        for (n637 = 0; n637 < 16; n637 = n637 + 1) 
        begin: outbit637
            assign data_11[n637 + d637*16 + c22*28*16] = data_11_array[c22][d637][n637];
        end
    endgenerate
    generate 
        localparam integer d638 = 22;
        for (n638 = 0; n638 < 16; n638 = n638 + 1) 
        begin: outbit638
            assign data_11[n638 + d638*16 + c22*28*16] = data_11_array[c22][d638][n638];
        end
    endgenerate
    generate 
        localparam integer d639 = 23;
        for (n639 = 0; n639 < 16; n639 = n639 + 1) 
        begin: outbit639
            assign data_11[n639 + d639*16 + c22*28*16] = data_11_array[c22][d639][n639];
        end
    endgenerate
    generate 
        localparam integer d640 = 24;
        for (n640 = 0; n640 < 16; n640 = n640 + 1) 
        begin: outbit640
            assign data_11[n640 + d640*16 + c22*28*16] = data_11_array[c22][d640][n640];
        end
    endgenerate
    generate 
        localparam integer d641 = 25;
        for (n641 = 0; n641 < 16; n641 = n641 + 1) 
        begin: outbit641
            assign data_11[n641 + d641*16 + c22*28*16] = data_11_array[c22][d641][n641];
        end
    endgenerate
    generate 
        localparam integer d642 = 26;
        for (n642 = 0; n642 < 16; n642 = n642 + 1) 
        begin: outbit642
            assign data_11[n642 + d642*16 + c22*28*16] = data_11_array[c22][d642][n642];
        end
    endgenerate
    generate 
        localparam integer d643 = 27;
        for (n643 = 0; n643 < 16; n643 = n643 + 1) 
        begin: outbit643
            assign data_11[n643 + d643*16 + c22*28*16] = data_11_array[c22][d643][n643];
        end
    endgenerate
    localparam integer c23 = 23;
    generate 
        localparam integer d644 = 0;
        for (n644 = 0; n644 < 16; n644 = n644 + 1) 
        begin: outbit644
            assign data_11[n644 + d644*16 + c23*28*16] = data_11_array[c23][d644][n644];
        end
    endgenerate
    generate 
        localparam integer d645 = 1;
        for (n645 = 0; n645 < 16; n645 = n645 + 1) 
        begin: outbit645
            assign data_11[n645 + d645*16 + c23*28*16] = data_11_array[c23][d645][n645];
        end
    endgenerate
    generate 
        localparam integer d646 = 2;
        for (n646 = 0; n646 < 16; n646 = n646 + 1) 
        begin: outbit646
            assign data_11[n646 + d646*16 + c23*28*16] = data_11_array[c23][d646][n646];
        end
    endgenerate
    generate 
        localparam integer d647 = 3;
        for (n647 = 0; n647 < 16; n647 = n647 + 1) 
        begin: outbit647
            assign data_11[n647 + d647*16 + c23*28*16] = data_11_array[c23][d647][n647];
        end
    endgenerate
    generate 
        localparam integer d648 = 4;
        for (n648 = 0; n648 < 16; n648 = n648 + 1) 
        begin: outbit648
            assign data_11[n648 + d648*16 + c23*28*16] = data_11_array[c23][d648][n648];
        end
    endgenerate
    generate 
        localparam integer d649 = 5;
        for (n649 = 0; n649 < 16; n649 = n649 + 1) 
        begin: outbit649
            assign data_11[n649 + d649*16 + c23*28*16] = data_11_array[c23][d649][n649];
        end
    endgenerate
    generate 
        localparam integer d650 = 6;
        for (n650 = 0; n650 < 16; n650 = n650 + 1) 
        begin: outbit650
            assign data_11[n650 + d650*16 + c23*28*16] = data_11_array[c23][d650][n650];
        end
    endgenerate
    generate 
        localparam integer d651 = 7;
        for (n651 = 0; n651 < 16; n651 = n651 + 1) 
        begin: outbit651
            assign data_11[n651 + d651*16 + c23*28*16] = data_11_array[c23][d651][n651];
        end
    endgenerate
    generate 
        localparam integer d652 = 8;
        for (n652 = 0; n652 < 16; n652 = n652 + 1) 
        begin: outbit652
            assign data_11[n652 + d652*16 + c23*28*16] = data_11_array[c23][d652][n652];
        end
    endgenerate
    generate 
        localparam integer d653 = 9;
        for (n653 = 0; n653 < 16; n653 = n653 + 1) 
        begin: outbit653
            assign data_11[n653 + d653*16 + c23*28*16] = data_11_array[c23][d653][n653];
        end
    endgenerate
    generate 
        localparam integer d654 = 10;
        for (n654 = 0; n654 < 16; n654 = n654 + 1) 
        begin: outbit654
            assign data_11[n654 + d654*16 + c23*28*16] = data_11_array[c23][d654][n654];
        end
    endgenerate
    generate 
        localparam integer d655 = 11;
        for (n655 = 0; n655 < 16; n655 = n655 + 1) 
        begin: outbit655
            assign data_11[n655 + d655*16 + c23*28*16] = data_11_array[c23][d655][n655];
        end
    endgenerate
    generate 
        localparam integer d656 = 12;
        for (n656 = 0; n656 < 16; n656 = n656 + 1) 
        begin: outbit656
            assign data_11[n656 + d656*16 + c23*28*16] = data_11_array[c23][d656][n656];
        end
    endgenerate
    generate 
        localparam integer d657 = 13;
        for (n657 = 0; n657 < 16; n657 = n657 + 1) 
        begin: outbit657
            assign data_11[n657 + d657*16 + c23*28*16] = data_11_array[c23][d657][n657];
        end
    endgenerate
    generate 
        localparam integer d658 = 14;
        for (n658 = 0; n658 < 16; n658 = n658 + 1) 
        begin: outbit658
            assign data_11[n658 + d658*16 + c23*28*16] = data_11_array[c23][d658][n658];
        end
    endgenerate
    generate 
        localparam integer d659 = 15;
        for (n659 = 0; n659 < 16; n659 = n659 + 1) 
        begin: outbit659
            assign data_11[n659 + d659*16 + c23*28*16] = data_11_array[c23][d659][n659];
        end
    endgenerate
    generate 
        localparam integer d660 = 16;
        for (n660 = 0; n660 < 16; n660 = n660 + 1) 
        begin: outbit660
            assign data_11[n660 + d660*16 + c23*28*16] = data_11_array[c23][d660][n660];
        end
    endgenerate
    generate 
        localparam integer d661 = 17;
        for (n661 = 0; n661 < 16; n661 = n661 + 1) 
        begin: outbit661
            assign data_11[n661 + d661*16 + c23*28*16] = data_11_array[c23][d661][n661];
        end
    endgenerate
    generate 
        localparam integer d662 = 18;
        for (n662 = 0; n662 < 16; n662 = n662 + 1) 
        begin: outbit662
            assign data_11[n662 + d662*16 + c23*28*16] = data_11_array[c23][d662][n662];
        end
    endgenerate
    generate 
        localparam integer d663 = 19;
        for (n663 = 0; n663 < 16; n663 = n663 + 1) 
        begin: outbit663
            assign data_11[n663 + d663*16 + c23*28*16] = data_11_array[c23][d663][n663];
        end
    endgenerate
    generate 
        localparam integer d664 = 20;
        for (n664 = 0; n664 < 16; n664 = n664 + 1) 
        begin: outbit664
            assign data_11[n664 + d664*16 + c23*28*16] = data_11_array[c23][d664][n664];
        end
    endgenerate
    generate 
        localparam integer d665 = 21;
        for (n665 = 0; n665 < 16; n665 = n665 + 1) 
        begin: outbit665
            assign data_11[n665 + d665*16 + c23*28*16] = data_11_array[c23][d665][n665];
        end
    endgenerate
    generate 
        localparam integer d666 = 22;
        for (n666 = 0; n666 < 16; n666 = n666 + 1) 
        begin: outbit666
            assign data_11[n666 + d666*16 + c23*28*16] = data_11_array[c23][d666][n666];
        end
    endgenerate
    generate 
        localparam integer d667 = 23;
        for (n667 = 0; n667 < 16; n667 = n667 + 1) 
        begin: outbit667
            assign data_11[n667 + d667*16 + c23*28*16] = data_11_array[c23][d667][n667];
        end
    endgenerate
    generate 
        localparam integer d668 = 24;
        for (n668 = 0; n668 < 16; n668 = n668 + 1) 
        begin: outbit668
            assign data_11[n668 + d668*16 + c23*28*16] = data_11_array[c23][d668][n668];
        end
    endgenerate
    generate 
        localparam integer d669 = 25;
        for (n669 = 0; n669 < 16; n669 = n669 + 1) 
        begin: outbit669
            assign data_11[n669 + d669*16 + c23*28*16] = data_11_array[c23][d669][n669];
        end
    endgenerate
    generate 
        localparam integer d670 = 26;
        for (n670 = 0; n670 < 16; n670 = n670 + 1) 
        begin: outbit670
            assign data_11[n670 + d670*16 + c23*28*16] = data_11_array[c23][d670][n670];
        end
    endgenerate
    generate 
        localparam integer d671 = 27;
        for (n671 = 0; n671 < 16; n671 = n671 + 1) 
        begin: outbit671
            assign data_11[n671 + d671*16 + c23*28*16] = data_11_array[c23][d671][n671];
        end
    endgenerate
    localparam integer c24 = 24;
    generate 
        localparam integer d672 = 0;
        for (n672 = 0; n672 < 16; n672 = n672 + 1) 
        begin: outbit672
            assign data_11[n672 + d672*16 + c24*28*16] = data_11_array[c24][d672][n672];
        end
    endgenerate
    generate 
        localparam integer d673 = 1;
        for (n673 = 0; n673 < 16; n673 = n673 + 1) 
        begin: outbit673
            assign data_11[n673 + d673*16 + c24*28*16] = data_11_array[c24][d673][n673];
        end
    endgenerate
    generate 
        localparam integer d674 = 2;
        for (n674 = 0; n674 < 16; n674 = n674 + 1) 
        begin: outbit674
            assign data_11[n674 + d674*16 + c24*28*16] = data_11_array[c24][d674][n674];
        end
    endgenerate
    generate 
        localparam integer d675 = 3;
        for (n675 = 0; n675 < 16; n675 = n675 + 1) 
        begin: outbit675
            assign data_11[n675 + d675*16 + c24*28*16] = data_11_array[c24][d675][n675];
        end
    endgenerate
    generate 
        localparam integer d676 = 4;
        for (n676 = 0; n676 < 16; n676 = n676 + 1) 
        begin: outbit676
            assign data_11[n676 + d676*16 + c24*28*16] = data_11_array[c24][d676][n676];
        end
    endgenerate
    generate 
        localparam integer d677 = 5;
        for (n677 = 0; n677 < 16; n677 = n677 + 1) 
        begin: outbit677
            assign data_11[n677 + d677*16 + c24*28*16] = data_11_array[c24][d677][n677];
        end
    endgenerate
    generate 
        localparam integer d678 = 6;
        for (n678 = 0; n678 < 16; n678 = n678 + 1) 
        begin: outbit678
            assign data_11[n678 + d678*16 + c24*28*16] = data_11_array[c24][d678][n678];
        end
    endgenerate
    generate 
        localparam integer d679 = 7;
        for (n679 = 0; n679 < 16; n679 = n679 + 1) 
        begin: outbit679
            assign data_11[n679 + d679*16 + c24*28*16] = data_11_array[c24][d679][n679];
        end
    endgenerate
    generate 
        localparam integer d680 = 8;
        for (n680 = 0; n680 < 16; n680 = n680 + 1) 
        begin: outbit680
            assign data_11[n680 + d680*16 + c24*28*16] = data_11_array[c24][d680][n680];
        end
    endgenerate
    generate 
        localparam integer d681 = 9;
        for (n681 = 0; n681 < 16; n681 = n681 + 1) 
        begin: outbit681
            assign data_11[n681 + d681*16 + c24*28*16] = data_11_array[c24][d681][n681];
        end
    endgenerate
    generate 
        localparam integer d682 = 10;
        for (n682 = 0; n682 < 16; n682 = n682 + 1) 
        begin: outbit682
            assign data_11[n682 + d682*16 + c24*28*16] = data_11_array[c24][d682][n682];
        end
    endgenerate
    generate 
        localparam integer d683 = 11;
        for (n683 = 0; n683 < 16; n683 = n683 + 1) 
        begin: outbit683
            assign data_11[n683 + d683*16 + c24*28*16] = data_11_array[c24][d683][n683];
        end
    endgenerate
    generate 
        localparam integer d684 = 12;
        for (n684 = 0; n684 < 16; n684 = n684 + 1) 
        begin: outbit684
            assign data_11[n684 + d684*16 + c24*28*16] = data_11_array[c24][d684][n684];
        end
    endgenerate
    generate 
        localparam integer d685 = 13;
        for (n685 = 0; n685 < 16; n685 = n685 + 1) 
        begin: outbit685
            assign data_11[n685 + d685*16 + c24*28*16] = data_11_array[c24][d685][n685];
        end
    endgenerate
    generate 
        localparam integer d686 = 14;
        for (n686 = 0; n686 < 16; n686 = n686 + 1) 
        begin: outbit686
            assign data_11[n686 + d686*16 + c24*28*16] = data_11_array[c24][d686][n686];
        end
    endgenerate
    generate 
        localparam integer d687 = 15;
        for (n687 = 0; n687 < 16; n687 = n687 + 1) 
        begin: outbit687
            assign data_11[n687 + d687*16 + c24*28*16] = data_11_array[c24][d687][n687];
        end
    endgenerate
    generate 
        localparam integer d688 = 16;
        for (n688 = 0; n688 < 16; n688 = n688 + 1) 
        begin: outbit688
            assign data_11[n688 + d688*16 + c24*28*16] = data_11_array[c24][d688][n688];
        end
    endgenerate
    generate 
        localparam integer d689 = 17;
        for (n689 = 0; n689 < 16; n689 = n689 + 1) 
        begin: outbit689
            assign data_11[n689 + d689*16 + c24*28*16] = data_11_array[c24][d689][n689];
        end
    endgenerate
    generate 
        localparam integer d690 = 18;
        for (n690 = 0; n690 < 16; n690 = n690 + 1) 
        begin: outbit690
            assign data_11[n690 + d690*16 + c24*28*16] = data_11_array[c24][d690][n690];
        end
    endgenerate
    generate 
        localparam integer d691 = 19;
        for (n691 = 0; n691 < 16; n691 = n691 + 1) 
        begin: outbit691
            assign data_11[n691 + d691*16 + c24*28*16] = data_11_array[c24][d691][n691];
        end
    endgenerate
    generate 
        localparam integer d692 = 20;
        for (n692 = 0; n692 < 16; n692 = n692 + 1) 
        begin: outbit692
            assign data_11[n692 + d692*16 + c24*28*16] = data_11_array[c24][d692][n692];
        end
    endgenerate
    generate 
        localparam integer d693 = 21;
        for (n693 = 0; n693 < 16; n693 = n693 + 1) 
        begin: outbit693
            assign data_11[n693 + d693*16 + c24*28*16] = data_11_array[c24][d693][n693];
        end
    endgenerate
    generate 
        localparam integer d694 = 22;
        for (n694 = 0; n694 < 16; n694 = n694 + 1) 
        begin: outbit694
            assign data_11[n694 + d694*16 + c24*28*16] = data_11_array[c24][d694][n694];
        end
    endgenerate
    generate 
        localparam integer d695 = 23;
        for (n695 = 0; n695 < 16; n695 = n695 + 1) 
        begin: outbit695
            assign data_11[n695 + d695*16 + c24*28*16] = data_11_array[c24][d695][n695];
        end
    endgenerate
    generate 
        localparam integer d696 = 24;
        for (n696 = 0; n696 < 16; n696 = n696 + 1) 
        begin: outbit696
            assign data_11[n696 + d696*16 + c24*28*16] = data_11_array[c24][d696][n696];
        end
    endgenerate
    generate 
        localparam integer d697 = 25;
        for (n697 = 0; n697 < 16; n697 = n697 + 1) 
        begin: outbit697
            assign data_11[n697 + d697*16 + c24*28*16] = data_11_array[c24][d697][n697];
        end
    endgenerate
    generate 
        localparam integer d698 = 26;
        for (n698 = 0; n698 < 16; n698 = n698 + 1) 
        begin: outbit698
            assign data_11[n698 + d698*16 + c24*28*16] = data_11_array[c24][d698][n698];
        end
    endgenerate
    generate 
        localparam integer d699 = 27;
        for (n699 = 0; n699 < 16; n699 = n699 + 1) 
        begin: outbit699
            assign data_11[n699 + d699*16 + c24*28*16] = data_11_array[c24][d699][n699];
        end
    endgenerate
    localparam integer c25 = 25;
    generate 
        localparam integer d700 = 0;
        for (n700 = 0; n700 < 16; n700 = n700 + 1) 
        begin: outbit700
            assign data_11[n700 + d700*16 + c25*28*16] = data_11_array[c25][d700][n700];
        end
    endgenerate
    generate 
        localparam integer d701 = 1;
        for (n701 = 0; n701 < 16; n701 = n701 + 1) 
        begin: outbit701
            assign data_11[n701 + d701*16 + c25*28*16] = data_11_array[c25][d701][n701];
        end
    endgenerate
    generate 
        localparam integer d702 = 2;
        for (n702 = 0; n702 < 16; n702 = n702 + 1) 
        begin: outbit702
            assign data_11[n702 + d702*16 + c25*28*16] = data_11_array[c25][d702][n702];
        end
    endgenerate
    generate 
        localparam integer d703 = 3;
        for (n703 = 0; n703 < 16; n703 = n703 + 1) 
        begin: outbit703
            assign data_11[n703 + d703*16 + c25*28*16] = data_11_array[c25][d703][n703];
        end
    endgenerate
    generate 
        localparam integer d704 = 4;
        for (n704 = 0; n704 < 16; n704 = n704 + 1) 
        begin: outbit704
            assign data_11[n704 + d704*16 + c25*28*16] = data_11_array[c25][d704][n704];
        end
    endgenerate
    generate 
        localparam integer d705 = 5;
        for (n705 = 0; n705 < 16; n705 = n705 + 1) 
        begin: outbit705
            assign data_11[n705 + d705*16 + c25*28*16] = data_11_array[c25][d705][n705];
        end
    endgenerate
    generate 
        localparam integer d706 = 6;
        for (n706 = 0; n706 < 16; n706 = n706 + 1) 
        begin: outbit706
            assign data_11[n706 + d706*16 + c25*28*16] = data_11_array[c25][d706][n706];
        end
    endgenerate
    generate 
        localparam integer d707 = 7;
        for (n707 = 0; n707 < 16; n707 = n707 + 1) 
        begin: outbit707
            assign data_11[n707 + d707*16 + c25*28*16] = data_11_array[c25][d707][n707];
        end
    endgenerate
    generate 
        localparam integer d708 = 8;
        for (n708 = 0; n708 < 16; n708 = n708 + 1) 
        begin: outbit708
            assign data_11[n708 + d708*16 + c25*28*16] = data_11_array[c25][d708][n708];
        end
    endgenerate
    generate 
        localparam integer d709 = 9;
        for (n709 = 0; n709 < 16; n709 = n709 + 1) 
        begin: outbit709
            assign data_11[n709 + d709*16 + c25*28*16] = data_11_array[c25][d709][n709];
        end
    endgenerate
    generate 
        localparam integer d710 = 10;
        for (n710 = 0; n710 < 16; n710 = n710 + 1) 
        begin: outbit710
            assign data_11[n710 + d710*16 + c25*28*16] = data_11_array[c25][d710][n710];
        end
    endgenerate
    generate 
        localparam integer d711 = 11;
        for (n711 = 0; n711 < 16; n711 = n711 + 1) 
        begin: outbit711
            assign data_11[n711 + d711*16 + c25*28*16] = data_11_array[c25][d711][n711];
        end
    endgenerate
    generate 
        localparam integer d712 = 12;
        for (n712 = 0; n712 < 16; n712 = n712 + 1) 
        begin: outbit712
            assign data_11[n712 + d712*16 + c25*28*16] = data_11_array[c25][d712][n712];
        end
    endgenerate
    generate 
        localparam integer d713 = 13;
        for (n713 = 0; n713 < 16; n713 = n713 + 1) 
        begin: outbit713
            assign data_11[n713 + d713*16 + c25*28*16] = data_11_array[c25][d713][n713];
        end
    endgenerate
    generate 
        localparam integer d714 = 14;
        for (n714 = 0; n714 < 16; n714 = n714 + 1) 
        begin: outbit714
            assign data_11[n714 + d714*16 + c25*28*16] = data_11_array[c25][d714][n714];
        end
    endgenerate
    generate 
        localparam integer d715 = 15;
        for (n715 = 0; n715 < 16; n715 = n715 + 1) 
        begin: outbit715
            assign data_11[n715 + d715*16 + c25*28*16] = data_11_array[c25][d715][n715];
        end
    endgenerate
    generate 
        localparam integer d716 = 16;
        for (n716 = 0; n716 < 16; n716 = n716 + 1) 
        begin: outbit716
            assign data_11[n716 + d716*16 + c25*28*16] = data_11_array[c25][d716][n716];
        end
    endgenerate
    generate 
        localparam integer d717 = 17;
        for (n717 = 0; n717 < 16; n717 = n717 + 1) 
        begin: outbit717
            assign data_11[n717 + d717*16 + c25*28*16] = data_11_array[c25][d717][n717];
        end
    endgenerate
    generate 
        localparam integer d718 = 18;
        for (n718 = 0; n718 < 16; n718 = n718 + 1) 
        begin: outbit718
            assign data_11[n718 + d718*16 + c25*28*16] = data_11_array[c25][d718][n718];
        end
    endgenerate
    generate 
        localparam integer d719 = 19;
        for (n719 = 0; n719 < 16; n719 = n719 + 1) 
        begin: outbit719
            assign data_11[n719 + d719*16 + c25*28*16] = data_11_array[c25][d719][n719];
        end
    endgenerate
    generate 
        localparam integer d720 = 20;
        for (n720 = 0; n720 < 16; n720 = n720 + 1) 
        begin: outbit720
            assign data_11[n720 + d720*16 + c25*28*16] = data_11_array[c25][d720][n720];
        end
    endgenerate
    generate 
        localparam integer d721 = 21;
        for (n721 = 0; n721 < 16; n721 = n721 + 1) 
        begin: outbit721
            assign data_11[n721 + d721*16 + c25*28*16] = data_11_array[c25][d721][n721];
        end
    endgenerate
    generate 
        localparam integer d722 = 22;
        for (n722 = 0; n722 < 16; n722 = n722 + 1) 
        begin: outbit722
            assign data_11[n722 + d722*16 + c25*28*16] = data_11_array[c25][d722][n722];
        end
    endgenerate
    generate 
        localparam integer d723 = 23;
        for (n723 = 0; n723 < 16; n723 = n723 + 1) 
        begin: outbit723
            assign data_11[n723 + d723*16 + c25*28*16] = data_11_array[c25][d723][n723];
        end
    endgenerate
    generate 
        localparam integer d724 = 24;
        for (n724 = 0; n724 < 16; n724 = n724 + 1) 
        begin: outbit724
            assign data_11[n724 + d724*16 + c25*28*16] = data_11_array[c25][d724][n724];
        end
    endgenerate
    generate 
        localparam integer d725 = 25;
        for (n725 = 0; n725 < 16; n725 = n725 + 1) 
        begin: outbit725
            assign data_11[n725 + d725*16 + c25*28*16] = data_11_array[c25][d725][n725];
        end
    endgenerate
    generate 
        localparam integer d726 = 26;
        for (n726 = 0; n726 < 16; n726 = n726 + 1) 
        begin: outbit726
            assign data_11[n726 + d726*16 + c25*28*16] = data_11_array[c25][d726][n726];
        end
    endgenerate
    generate 
        localparam integer d727 = 27;
        for (n727 = 0; n727 < 16; n727 = n727 + 1) 
        begin: outbit727
            assign data_11[n727 + d727*16 + c25*28*16] = data_11_array[c25][d727][n727];
        end
    endgenerate
    localparam integer c26 = 26;
    generate 
        localparam integer d728 = 0;
        for (n728 = 0; n728 < 16; n728 = n728 + 1) 
        begin: outbit728
            assign data_11[n728 + d728*16 + c26*28*16] = data_11_array[c26][d728][n728];
        end
    endgenerate
    generate 
        localparam integer d729 = 1;
        for (n729 = 0; n729 < 16; n729 = n729 + 1) 
        begin: outbit729
            assign data_11[n729 + d729*16 + c26*28*16] = data_11_array[c26][d729][n729];
        end
    endgenerate
    generate 
        localparam integer d730 = 2;
        for (n730 = 0; n730 < 16; n730 = n730 + 1) 
        begin: outbit730
            assign data_11[n730 + d730*16 + c26*28*16] = data_11_array[c26][d730][n730];
        end
    endgenerate
    generate 
        localparam integer d731 = 3;
        for (n731 = 0; n731 < 16; n731 = n731 + 1) 
        begin: outbit731
            assign data_11[n731 + d731*16 + c26*28*16] = data_11_array[c26][d731][n731];
        end
    endgenerate
    generate 
        localparam integer d732 = 4;
        for (n732 = 0; n732 < 16; n732 = n732 + 1) 
        begin: outbit732
            assign data_11[n732 + d732*16 + c26*28*16] = data_11_array[c26][d732][n732];
        end
    endgenerate
    generate 
        localparam integer d733 = 5;
        for (n733 = 0; n733 < 16; n733 = n733 + 1) 
        begin: outbit733
            assign data_11[n733 + d733*16 + c26*28*16] = data_11_array[c26][d733][n733];
        end
    endgenerate
    generate 
        localparam integer d734 = 6;
        for (n734 = 0; n734 < 16; n734 = n734 + 1) 
        begin: outbit734
            assign data_11[n734 + d734*16 + c26*28*16] = data_11_array[c26][d734][n734];
        end
    endgenerate
    generate 
        localparam integer d735 = 7;
        for (n735 = 0; n735 < 16; n735 = n735 + 1) 
        begin: outbit735
            assign data_11[n735 + d735*16 + c26*28*16] = data_11_array[c26][d735][n735];
        end
    endgenerate
    generate 
        localparam integer d736 = 8;
        for (n736 = 0; n736 < 16; n736 = n736 + 1) 
        begin: outbit736
            assign data_11[n736 + d736*16 + c26*28*16] = data_11_array[c26][d736][n736];
        end
    endgenerate
    generate 
        localparam integer d737 = 9;
        for (n737 = 0; n737 < 16; n737 = n737 + 1) 
        begin: outbit737
            assign data_11[n737 + d737*16 + c26*28*16] = data_11_array[c26][d737][n737];
        end
    endgenerate
    generate 
        localparam integer d738 = 10;
        for (n738 = 0; n738 < 16; n738 = n738 + 1) 
        begin: outbit738
            assign data_11[n738 + d738*16 + c26*28*16] = data_11_array[c26][d738][n738];
        end
    endgenerate
    generate 
        localparam integer d739 = 11;
        for (n739 = 0; n739 < 16; n739 = n739 + 1) 
        begin: outbit739
            assign data_11[n739 + d739*16 + c26*28*16] = data_11_array[c26][d739][n739];
        end
    endgenerate
    generate 
        localparam integer d740 = 12;
        for (n740 = 0; n740 < 16; n740 = n740 + 1) 
        begin: outbit740
            assign data_11[n740 + d740*16 + c26*28*16] = data_11_array[c26][d740][n740];
        end
    endgenerate
    generate 
        localparam integer d741 = 13;
        for (n741 = 0; n741 < 16; n741 = n741 + 1) 
        begin: outbit741
            assign data_11[n741 + d741*16 + c26*28*16] = data_11_array[c26][d741][n741];
        end
    endgenerate
    generate 
        localparam integer d742 = 14;
        for (n742 = 0; n742 < 16; n742 = n742 + 1) 
        begin: outbit742
            assign data_11[n742 + d742*16 + c26*28*16] = data_11_array[c26][d742][n742];
        end
    endgenerate
    generate 
        localparam integer d743 = 15;
        for (n743 = 0; n743 < 16; n743 = n743 + 1) 
        begin: outbit743
            assign data_11[n743 + d743*16 + c26*28*16] = data_11_array[c26][d743][n743];
        end
    endgenerate
    generate 
        localparam integer d744 = 16;
        for (n744 = 0; n744 < 16; n744 = n744 + 1) 
        begin: outbit744
            assign data_11[n744 + d744*16 + c26*28*16] = data_11_array[c26][d744][n744];
        end
    endgenerate
    generate 
        localparam integer d745 = 17;
        for (n745 = 0; n745 < 16; n745 = n745 + 1) 
        begin: outbit745
            assign data_11[n745 + d745*16 + c26*28*16] = data_11_array[c26][d745][n745];
        end
    endgenerate
    generate 
        localparam integer d746 = 18;
        for (n746 = 0; n746 < 16; n746 = n746 + 1) 
        begin: outbit746
            assign data_11[n746 + d746*16 + c26*28*16] = data_11_array[c26][d746][n746];
        end
    endgenerate
    generate 
        localparam integer d747 = 19;
        for (n747 = 0; n747 < 16; n747 = n747 + 1) 
        begin: outbit747
            assign data_11[n747 + d747*16 + c26*28*16] = data_11_array[c26][d747][n747];
        end
    endgenerate
    generate 
        localparam integer d748 = 20;
        for (n748 = 0; n748 < 16; n748 = n748 + 1) 
        begin: outbit748
            assign data_11[n748 + d748*16 + c26*28*16] = data_11_array[c26][d748][n748];
        end
    endgenerate
    generate 
        localparam integer d749 = 21;
        for (n749 = 0; n749 < 16; n749 = n749 + 1) 
        begin: outbit749
            assign data_11[n749 + d749*16 + c26*28*16] = data_11_array[c26][d749][n749];
        end
    endgenerate
    generate 
        localparam integer d750 = 22;
        for (n750 = 0; n750 < 16; n750 = n750 + 1) 
        begin: outbit750
            assign data_11[n750 + d750*16 + c26*28*16] = data_11_array[c26][d750][n750];
        end
    endgenerate
    generate 
        localparam integer d751 = 23;
        for (n751 = 0; n751 < 16; n751 = n751 + 1) 
        begin: outbit751
            assign data_11[n751 + d751*16 + c26*28*16] = data_11_array[c26][d751][n751];
        end
    endgenerate
    generate 
        localparam integer d752 = 24;
        for (n752 = 0; n752 < 16; n752 = n752 + 1) 
        begin: outbit752
            assign data_11[n752 + d752*16 + c26*28*16] = data_11_array[c26][d752][n752];
        end
    endgenerate
    generate 
        localparam integer d753 = 25;
        for (n753 = 0; n753 < 16; n753 = n753 + 1) 
        begin: outbit753
            assign data_11[n753 + d753*16 + c26*28*16] = data_11_array[c26][d753][n753];
        end
    endgenerate
    generate 
        localparam integer d754 = 26;
        for (n754 = 0; n754 < 16; n754 = n754 + 1) 
        begin: outbit754
            assign data_11[n754 + d754*16 + c26*28*16] = data_11_array[c26][d754][n754];
        end
    endgenerate
    generate 
        localparam integer d755 = 27;
        for (n755 = 0; n755 < 16; n755 = n755 + 1) 
        begin: outbit755
            assign data_11[n755 + d755*16 + c26*28*16] = data_11_array[c26][d755][n755];
        end
    endgenerate
    localparam integer c27 = 27;
    generate 
        localparam integer d756 = 0;
        for (n756 = 0; n756 < 16; n756 = n756 + 1) 
        begin: outbit756
            assign data_11[n756 + d756*16 + c27*28*16] = data_11_array[c27][d756][n756];
        end
    endgenerate
    generate 
        localparam integer d757 = 1;
        for (n757 = 0; n757 < 16; n757 = n757 + 1) 
        begin: outbit757
            assign data_11[n757 + d757*16 + c27*28*16] = data_11_array[c27][d757][n757];
        end
    endgenerate
    generate 
        localparam integer d758 = 2;
        for (n758 = 0; n758 < 16; n758 = n758 + 1) 
        begin: outbit758
            assign data_11[n758 + d758*16 + c27*28*16] = data_11_array[c27][d758][n758];
        end
    endgenerate
    generate 
        localparam integer d759 = 3;
        for (n759 = 0; n759 < 16; n759 = n759 + 1) 
        begin: outbit759
            assign data_11[n759 + d759*16 + c27*28*16] = data_11_array[c27][d759][n759];
        end
    endgenerate
    generate 
        localparam integer d760 = 4;
        for (n760 = 0; n760 < 16; n760 = n760 + 1) 
        begin: outbit760
            assign data_11[n760 + d760*16 + c27*28*16] = data_11_array[c27][d760][n760];
        end
    endgenerate
    generate 
        localparam integer d761 = 5;
        for (n761 = 0; n761 < 16; n761 = n761 + 1) 
        begin: outbit761
            assign data_11[n761 + d761*16 + c27*28*16] = data_11_array[c27][d761][n761];
        end
    endgenerate
    generate 
        localparam integer d762 = 6;
        for (n762 = 0; n762 < 16; n762 = n762 + 1) 
        begin: outbit762
            assign data_11[n762 + d762*16 + c27*28*16] = data_11_array[c27][d762][n762];
        end
    endgenerate
    generate 
        localparam integer d763 = 7;
        for (n763 = 0; n763 < 16; n763 = n763 + 1) 
        begin: outbit763
            assign data_11[n763 + d763*16 + c27*28*16] = data_11_array[c27][d763][n763];
        end
    endgenerate
    generate 
        localparam integer d764 = 8;
        for (n764 = 0; n764 < 16; n764 = n764 + 1) 
        begin: outbit764
            assign data_11[n764 + d764*16 + c27*28*16] = data_11_array[c27][d764][n764];
        end
    endgenerate
    generate 
        localparam integer d765 = 9;
        for (n765 = 0; n765 < 16; n765 = n765 + 1) 
        begin: outbit765
            assign data_11[n765 + d765*16 + c27*28*16] = data_11_array[c27][d765][n765];
        end
    endgenerate
    generate 
        localparam integer d766 = 10;
        for (n766 = 0; n766 < 16; n766 = n766 + 1) 
        begin: outbit766
            assign data_11[n766 + d766*16 + c27*28*16] = data_11_array[c27][d766][n766];
        end
    endgenerate
    generate 
        localparam integer d767 = 11;
        for (n767 = 0; n767 < 16; n767 = n767 + 1) 
        begin: outbit767
            assign data_11[n767 + d767*16 + c27*28*16] = data_11_array[c27][d767][n767];
        end
    endgenerate
    generate 
        localparam integer d768 = 12;
        for (n768 = 0; n768 < 16; n768 = n768 + 1) 
        begin: outbit768
            assign data_11[n768 + d768*16 + c27*28*16] = data_11_array[c27][d768][n768];
        end
    endgenerate
    generate 
        localparam integer d769 = 13;
        for (n769 = 0; n769 < 16; n769 = n769 + 1) 
        begin: outbit769
            assign data_11[n769 + d769*16 + c27*28*16] = data_11_array[c27][d769][n769];
        end
    endgenerate
    generate 
        localparam integer d770 = 14;
        for (n770 = 0; n770 < 16; n770 = n770 + 1) 
        begin: outbit770
            assign data_11[n770 + d770*16 + c27*28*16] = data_11_array[c27][d770][n770];
        end
    endgenerate
    generate 
        localparam integer d771 = 15;
        for (n771 = 0; n771 < 16; n771 = n771 + 1) 
        begin: outbit771
            assign data_11[n771 + d771*16 + c27*28*16] = data_11_array[c27][d771][n771];
        end
    endgenerate
    generate 
        localparam integer d772 = 16;
        for (n772 = 0; n772 < 16; n772 = n772 + 1) 
        begin: outbit772
            assign data_11[n772 + d772*16 + c27*28*16] = data_11_array[c27][d772][n772];
        end
    endgenerate
    generate 
        localparam integer d773 = 17;
        for (n773 = 0; n773 < 16; n773 = n773 + 1) 
        begin: outbit773
            assign data_11[n773 + d773*16 + c27*28*16] = data_11_array[c27][d773][n773];
        end
    endgenerate
    generate 
        localparam integer d774 = 18;
        for (n774 = 0; n774 < 16; n774 = n774 + 1) 
        begin: outbit774
            assign data_11[n774 + d774*16 + c27*28*16] = data_11_array[c27][d774][n774];
        end
    endgenerate
    generate 
        localparam integer d775 = 19;
        for (n775 = 0; n775 < 16; n775 = n775 + 1) 
        begin: outbit775
            assign data_11[n775 + d775*16 + c27*28*16] = data_11_array[c27][d775][n775];
        end
    endgenerate
    generate 
        localparam integer d776 = 20;
        for (n776 = 0; n776 < 16; n776 = n776 + 1) 
        begin: outbit776
            assign data_11[n776 + d776*16 + c27*28*16] = data_11_array[c27][d776][n776];
        end
    endgenerate
    generate 
        localparam integer d777 = 21;
        for (n777 = 0; n777 < 16; n777 = n777 + 1) 
        begin: outbit777
            assign data_11[n777 + d777*16 + c27*28*16] = data_11_array[c27][d777][n777];
        end
    endgenerate
    generate 
        localparam integer d778 = 22;
        for (n778 = 0; n778 < 16; n778 = n778 + 1) 
        begin: outbit778
            assign data_11[n778 + d778*16 + c27*28*16] = data_11_array[c27][d778][n778];
        end
    endgenerate
    generate 
        localparam integer d779 = 23;
        for (n779 = 0; n779 < 16; n779 = n779 + 1) 
        begin: outbit779
            assign data_11[n779 + d779*16 + c27*28*16] = data_11_array[c27][d779][n779];
        end
    endgenerate
    generate 
        localparam integer d780 = 24;
        for (n780 = 0; n780 < 16; n780 = n780 + 1) 
        begin: outbit780
            assign data_11[n780 + d780*16 + c27*28*16] = data_11_array[c27][d780][n780];
        end
    endgenerate
    generate 
        localparam integer d781 = 25;
        for (n781 = 0; n781 < 16; n781 = n781 + 1) 
        begin: outbit781
            assign data_11[n781 + d781*16 + c27*28*16] = data_11_array[c27][d781][n781];
        end
    endgenerate
    generate 
        localparam integer d782 = 26;
        for (n782 = 0; n782 < 16; n782 = n782 + 1) 
        begin: outbit782
            assign data_11[n782 + d782*16 + c27*28*16] = data_11_array[c27][d782][n782];
        end
    endgenerate
    generate 
        localparam integer d783 = 27;
        for (n783 = 0; n783 < 16; n783 = n783 + 1) 
        begin: outbit783
            assign data_11[n783 + d783*16 + c27*28*16] = data_11_array[c27][d783][n783];
        end
    endgenerate

 
endmodule

////CONVOLUTION LAYER 1 | FEATURE MAP 3
module Conv1_feature3 (
    data,
    feature3Weight_0,
    feature3Weight_1,
    feature3Weight_2,
    feature3Weight_3,
    feature3Weight_4,
    feature3Weight_5,
    feature3Weight_6,
    feature3Weight_7,
    feature3Weight_8,
    feature3Weight_9,
    feature3Weight_10,
    feature3Weight_11,
    feature3Weight_12,
    feature3Weight_13,
    feature3Weight_14,
    feature3Weight_15,
    feature3Weight_16,
    feature3Weight_17,
    feature3Weight_18,
    feature3Weight_19,
    feature3Weight_20,
    feature3Weight_21,
    feature3Weight_22,
    feature3Weight_23,
    feature3Weight_24,
    feature3Bias,
    data_11);

  parameter TEST_DATA = 784*16,
    FP_LENGTH = 16;
  input [TEST_DATA - 1:0] data;
  input [FP_LENGTH - 1:0] feature3Weight_0, feature3Weight_1, feature3Weight_2, feature3Weight_3, feature3Weight_4, feature3Weight_5, feature3Weight_6, feature3Weight_7, feature3Weight_8, feature3Weight_9, feature3Weight_10, feature3Weight_11, feature3Weight_12, feature3Weight_13, feature3Weight_14, feature3Weight_15, feature3Weight_16, feature3Weight_17, feature3Weight_18, feature3Weight_19, feature3Weight_20, feature3Weight_21, feature3Weight_22, feature3Weight_23, feature3Weight_24, feature3Bias;
  output [576*16 - 1:0] data_11;    
  
  wire [FP_LENGTH - 1:0] data_array [0:27][0:27];
  wire [FP_LENGTH - 1:0] data_11_array [0:23][0:23];
  wire [FP_LENGTH - 1:0] multi0 [0:24][0:23], multi1 [0:24][0:23], multi2 [0:24][0:23], multi3 [0:24][0:23], multi4 [0:24][0:23], multi5 [0:24][0:23], multi6 [0:24][0:23], multi7 [0:24][0:23], multi8 [0:24][0:23], multi9 [0:24][0:23], multi10 [0:24][0:23], multi11 [0:24][0:23], multi12 [0:24][0:23], multi13 [0:24][0:23], multi14 [0:24][0:23], multi15 [0:24][0:23], multi16 [0:24][0:23], multi17 [0:24][0:23], multi18 [0:24][0:23], multi19 [0:24][0:23], multi20 [0:24][0:23], multi21 [0:24][0:23], multi22 [0:24][0:23], multi23 [0:24][0:23], multi24 [0:24][0:23];
  wire [FP_LENGTH - 1:0] sum0 [0:23][0:23], sum1 [0:23][0:23], sum2 [0:23][0:23], sum3 [0:23][0:23], sum4 [0:23][0:23], sum5 [0:23][0:23], sum6 [0:23][0:23], sum7 [0:23][0:23], sum8 [0:23][0:23], sum9 [0:23][0:23], sum10 [0:23][0:23], sum11 [0:23][0:23], sum12 [0:23][0:23], sum13 [0:23][0:23], sum14 [0:23][0:23], sum15 [0:23][0:23], sum16 [0:23][0:23], sum17 [0:23][0:23], sum18 [0:23][0:23], sum19 [0:23][0:23], sum20 [0:23][0:23], sum21 [0:23][0:23], sum22 [0:23][0:23], sum23 [0:23][0:23], sum24 [0:23][0:23];
//  integer a, b, c; ///a = ROW, b = COLUMN, c = 16 bit Value
  
//  initial begin
//    for (a = 0; a < 28; a = a + 1) begin
//        for (b = 0; b < 28; b = b + 1) begin
//            for (c = 15; c >= 0; c = c - 1) begin
//                data_array[a][b][c] = data[c + b*16 + a*28*16];
//            end
//        end
//    end
    
//    forever begin
//        for (a = 0; a < 28; a = a + 1) begin
//            for (b = 0; b < 28; b = b + 1) begin
//                for (c = 15; c >= 0; c = c - 1) begin
//                   data_11[c + b*16 + a*28*16] = data_11_array[a][b][c];
//                end
//            end
//        end
//    end
//  end
  
  
  
genvar i0, i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21, i22, i23, m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15,m16,m17,m18,m19,m20,m21,m22,m23,m24,m25,m26,m27,m28,m29,m30,m31,m32,m33,m34,m35,m36,m37,m38,m39,m40,m41,m42,m43,m44,m45,m46,m47,m48,m49,m50,m51,m52,m53,m54,m55,m56,m57,m58,m59,m60,m61,m62,m63,m64,m65,m66,m67,m68,m69,m70,m71,m72,m73,m74,m75,m76,m77,m78,m79,m80,m81,m82,m83,m84,m85,m86,m87,m88,m89,m90,m91,m92,m93,m94,m95,m96,m97,m98,m99,m100,m101,m102,m103,m104,m105,m106,m107,m108,m109,m110,m111,m112,m113,m114,m115,m116,m117,m118,m119,m120,m121,m122,m123,m124,m125,m126,m127,m128,m129,m130,m131,m132,m133,m134,m135,m136,m137,m138,m139,m140,m141,m142,m143,m144,m145,m146,m147,m148,m149,m150,m151,m152,m153,m154,m155,m156,m157,m158,m159,m160,m161,m162,m163,m164,m165,m166,m167,m168,m169,m170,m171,m172,m173,m174,m175,m176,m177,m178,m179,m180,m181,m182,m183,m184,m185,m186,m187,m188,m189,m190,m191,m192,m193,m194,m195,m196,m197,m198,m199,m200,m201,m202,m203,m204,m205,m206,m207,m208,m209,m210,m211,m212,m213,m214,m215,m216,m217,m218,m219,m220,m221,m222,m223,m224,m225,m226,m227,m228,m229,m230,m231,m232,m233,m234,m235,m236,m237,m238,m239,m240,m241,m242,m243,m244,m245,m246,m247,m248,m249,m250,m251,m252,m253,m254,m255,m256,m257,m258,m259,m260,m261,m262,m263,m264,m265,m266,m267,m268,m269,m270,m271,m272,m273,m274,m275,m276,m277,m278,m279,m280,m281,m282,m283,m284,m285,m286,m287,m288,m289,m290,m291,m292,m293,m294,m295,m296,m297,m298,m299,m300,m301,m302,m303,m304,m305,m306,m307,m308,m309,m310,m311,m312,m313,m314,m315,m316,m317,m318,m319,m320,m321,m322,m323,m324,m325,m326,m327,m328,m329,m330,m331,m332,m333,m334,m335,m336,m337,m338,m339,m340,m341,m342,m343,m344,m345,m346,m347,m348,m349,m350,m351,m352,m353,m354,m355,m356,m357,m358,m359,m360,m361,m362,m363,m364,m365,m366,m367,m368,m369,m370,m371,m372,m373,m374,m375,m376,m377,m378,m379,m380,m381,m382,m383,m384,m385,m386,m387,m388,m389,m390,m391,m392,m393,m394,m395,m396,m397,m398,m399,m400,m401,m402,m403,m404,m405,m406,m407,m408,m409,m410,m411,m412,m413,m414,m415,m416,m417,m418,m419,m420,m421,m422,m423,m424,m425,m426,m427,m428,m429,m430,m431,m432,m433,m434,m435,m436,m437,m438,m439,m440,m441,m442,m443,m444,m445,m446,m447,m448,m449,m450,m451,m452,m453,m454,m455,m456,m457,m458,m459,m460,m461,m462,m463,m464,m465,m466,m467,m468,m469,m470,m471,m472,m473,m474,m475,m476,m477,m478,m479,m480,m481,m482,m483,m484,m485,m486,m487,m488,m489,m490,m491,m492,m493,m494,m495,m496,m497,m498,m499,m500,m501,m502,m503,m504,m505,m506,m507,m508,m509,m510,m511,m512,m513,m514,m515,m516,m517,m518,m519,m520,m521,m522,m523,m524,m525,m526,m527,m528,m529,m530,m531,m532,m533,m534,m535,m536,m537,m538,m539,m540,m541,m542,m543,m544,m545,m546,m547,m548,m549,m550,m551,m552,m553,m554,m555,m556,m557,m558,m559,m560,m561,m562,m563,m564,m565,m566,m567,m568,m569,m570,m571,m572,m573,m574,m575,m576,m577,m578,m579,m580,m581,m582,m583,m584,m585,m586,m587,m588,m589,m590,m591,m592,m593,m594,m595,m596,m597,m598,m599,m600,m601,m602,m603,m604,m605,m606,m607,m608,m609,m610,m611,m612,m613,m614,m615,m616,m617,m618,m619,m620,m621,m622,m623,m624,m625,m626,m627,m628,m629,m630,m631,m632,m633,m634,m635,m636,m637,m638,m639,m640,m641,m642,m643,m644,m645,m646,m647,m648,m649,m650,m651,m652,m653,m654,m655,m656,m657,m658,m659,m660,m661,m662,m663,m664,m665,m666,m667,m668,m669,m670,m671,m672,m673,m674,m675,m676,m677,m678,m679,m680,m681,m682,m683,m684,m685,m686,m687,m688,m689,m690,m691,m692,m693,m694,m695,m696,m697,m698,m699,m700,m701,m702,m703,m704,m705,m706,m707,m708,m709,m710,m711,m712,m713,m714,m715,m716,m717,m718,m719,m720,m721,m722,m723,m724,m725,m726,m727,m728,m729,m730,m731,m732,m733,m734,m735,m736,m737,m738,m739,m740,m741,m742,m743,m744,m745,m746,m747,m748,m749,m750,m751,m752,m753,m754,m755,m756,m757,m758,m759,m760,m761,m762,m763,m764,m765,m766,m767,m768,m769,m770,m771,m772,m773,m774,m775,m776,m777,m778,m779,m780,m781,m782,m783,n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n50,n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80,n81,n82,n83,n84,n85,n86,n87,n88,n89,n90,n91,n92,n93,n94,n95,n96,n97,n98,n99,n100,n101,n102,n103,n104,n105,n106,n107,n108,n109,n110,n111,n112,n113,n114,n115,n116,n117,n118,n119,n120,n121,n122,n123,n124,n125,n126,n127,n128,n129,n130,n131,n132,n133,n134,n135,n136,n137,n138,n139,n140,n141,n142,n143,n144,n145,n146,n147,n148,n149,n150,n151,n152,n153,n154,n155,n156,n157,n158,n159,n160,n161,n162,n163,n164,n165,n166,n167,n168,n169,n170,n171,n172,n173,n174,n175,n176,n177,n178,n179,n180,n181,n182,n183,n184,n185,n186,n187,n188,n189,n190,n191,n192,n193,n194,n195,n196,n197,n198,n199,n200,n201,n202,n203,n204,n205,n206,n207,n208,n209,n210,n211,n212,n213,n214,n215,n216,n217,n218,n219,n220,n221,n222,n223,n224,n225,n226,n227,n228,n229,n230,n231,n232,n233,n234,n235,n236,n237,n238,n239,n240,n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,n251,n252,n253,n254,n255,n256,n257,n258,n259,n260,n261,n262,n263,n264,n265,n266,n267,n268,n269,n270,n271,n272,n273,n274,n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,n330,n331,n332,n333,n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,n345,n346,n347,n348,n349,n350,n351,n352,n353,n354,n355,n356,n357,n358,n359,n360,n361,n362,n363,n364,n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,n385,n386,n387,n388,n389,n390,n391,n392,n393,n394,n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,n415,n416,n417,n418,n419,n420,n421,n422,n423,n424,n425,n426,n427,n428,n429,n430,n431,n432,n433,n434,n435,n436,n437,n438,n439,n440,n441,n442,n443,n444,n445,n446,n447,n448,n449,n450,n451,n452,n453,n454,n455,n456,n457,n458,n459,n460,n461,n462,n463,n464,n465,n466,n467,n468,n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,n479,n480,n481,n482,n483,n484,n485,n486,n487,n488,n489,n490,n491,n492,n493,n494,n495,n496,n497,n498,n499,n500,n501,n502,n503,n504,n505,n506,n507,n508,n509,n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,n559,n560,n561,n562,n563,n564,n565,n566,n567,n568,n569,n570,n571,n572,n573,n574,n575,n576,n577,n578,n579,n580,n581,n582,n583,n584,n585,n586,n587,n588,n589,n590,n591,n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,n612,n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,n623,n624,n625,n626,n627,n628,n629,n630,n631,n632,n633,n634,n635,n636,n637,n638,n639,n640,n641,n642,n643,n644,n645,n646,n647,n648,n649,n650,n651,n652,n653,n654,n655,n656,n657,n658,n659,n660,n661,n662,n663,n664,n665,n666,n667,n668,n669,n670,n671,n672,n673,n674,n675,n676,n677,n678,n679,n680,n681,n682,n683,n684,n685,n686,n687,n688,n689,n690,n691,n692,n693,n694,n695,n696,n697,n698,n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,n709,n710,n711,n712,n713,n714,n715,n716,n717,n718,n719,n720,n721,n722,n723,n724,n725,n726,n727,n728,n729,n730,n731,n732,n733,n734,n735,n736,n737,n738,n739,n740,n741,n742,n743,n744,n745,n746,n747,n748,n749,n750,n751,n752,n753,n754,n755,n756,n757,n758,n759,n760,n761,n762,n763,n764,n765,n766,n767,n768,n769,n770,n771,n772,n773,n774,n775,n776,n777,n778,n779,n780,n781,n782,n783;
  
  localparam integer a0 = 0;
    generate 
        localparam integer b0 = 0;
        for (m0 = 0; m0 < 16; m0 = m0 + 1) 
        begin: inbit0
            assign data_11[m0 + b0*16 + a0*28*16] = data_11_array[a0][b0][m0];
        end
    endgenerate
    generate 
        localparam integer b1 = 1;
        for (m1 = 0; m1 < 16; m1 = m1 + 1) 
        begin: inbit1
            assign data_11[m1 + b1*16 + a0*28*16] = data_11_array[a0][b1][m1];
        end
    endgenerate
    generate 
        localparam integer b2 = 2;
        for (m2 = 0; m2 < 16; m2 = m2 + 1) 
        begin: inbit2
            assign data_11[m2 + b2*16 + a0*28*16] = data_11_array[a0][b2][m2];
        end
    endgenerate
    generate 
        localparam integer b3 = 3;
        for (m3 = 0; m3 < 16; m3 = m3 + 1) 
        begin: inbit3
            assign data_11[m3 + b3*16 + a0*28*16] = data_11_array[a0][b3][m3];
        end
    endgenerate
    generate 
        localparam integer b4 = 4;
        for (m4 = 0; m4 < 16; m4 = m4 + 1) 
        begin: inbit4
            assign data_11[m4 + b4*16 + a0*28*16] = data_11_array[a0][b4][m4];
        end
    endgenerate
    generate 
        localparam integer b5 = 5;
        for (m5 = 0; m5 < 16; m5 = m5 + 1) 
        begin: inbit5
            assign data_11[m5 + b5*16 + a0*28*16] = data_11_array[a0][b5][m5];
        end
    endgenerate
    generate 
        localparam integer b6 = 6;
        for (m6 = 0; m6 < 16; m6 = m6 + 1) 
        begin: inbit6
            assign data_11[m6 + b6*16 + a0*28*16] = data_11_array[a0][b6][m6];
        end
    endgenerate
    generate 
        localparam integer b7 = 7;
        for (m7 = 0; m7 < 16; m7 = m7 + 1) 
        begin: inbit7
            assign data_11[m7 + b7*16 + a0*28*16] = data_11_array[a0][b7][m7];
        end
    endgenerate
    generate 
        localparam integer b8 = 8;
        for (m8 = 0; m8 < 16; m8 = m8 + 1) 
        begin: inbit8
            assign data_11[m8 + b8*16 + a0*28*16] = data_11_array[a0][b8][m8];
        end
    endgenerate
    generate 
        localparam integer b9 = 9;
        for (m9 = 0; m9 < 16; m9 = m9 + 1) 
        begin: inbit9
            assign data_11[m9 + b9*16 + a0*28*16] = data_11_array[a0][b9][m9];
        end
    endgenerate
    generate 
        localparam integer b10 = 10;
        for (m10 = 0; m10 < 16; m10 = m10 + 1) 
        begin: inbit10
            assign data_11[m10 + b10*16 + a0*28*16] = data_11_array[a0][b10][m10];
        end
    endgenerate
    generate 
        localparam integer b11 = 11;
        for (m11 = 0; m11 < 16; m11 = m11 + 1) 
        begin: inbit11
            assign data_11[m11 + b11*16 + a0*28*16] = data_11_array[a0][b11][m11];
        end
    endgenerate
    generate 
        localparam integer b12 = 12;
        for (m12 = 0; m12 < 16; m12 = m12 + 1) 
        begin: inbit12
            assign data_11[m12 + b12*16 + a0*28*16] = data_11_array[a0][b12][m12];
        end
    endgenerate
    generate 
        localparam integer b13 = 13;
        for (m13 = 0; m13 < 16; m13 = m13 + 1) 
        begin: inbit13
            assign data_11[m13 + b13*16 + a0*28*16] = data_11_array[a0][b13][m13];
        end
    endgenerate
    generate 
        localparam integer b14 = 14;
        for (m14 = 0; m14 < 16; m14 = m14 + 1) 
        begin: inbit14
            assign data_11[m14 + b14*16 + a0*28*16] = data_11_array[a0][b14][m14];
        end
    endgenerate
    generate 
        localparam integer b15 = 15;
        for (m15 = 0; m15 < 16; m15 = m15 + 1) 
        begin: inbit15
            assign data_11[m15 + b15*16 + a0*28*16] = data_11_array[a0][b15][m15];
        end
    endgenerate
    generate 
        localparam integer b16 = 16;
        for (m16 = 0; m16 < 16; m16 = m16 + 1) 
        begin: inbit16
            assign data_11[m16 + b16*16 + a0*28*16] = data_11_array[a0][b16][m16];
        end
    endgenerate
    generate 
        localparam integer b17 = 17;
        for (m17 = 0; m17 < 16; m17 = m17 + 1) 
        begin: inbit17
            assign data_11[m17 + b17*16 + a0*28*16] = data_11_array[a0][b17][m17];
        end
    endgenerate
    generate 
        localparam integer b18 = 18;
        for (m18 = 0; m18 < 16; m18 = m18 + 1) 
        begin: inbit18
            assign data_11[m18 + b18*16 + a0*28*16] = data_11_array[a0][b18][m18];
        end
    endgenerate
    generate 
        localparam integer b19 = 19;
        for (m19 = 0; m19 < 16; m19 = m19 + 1) 
        begin: inbit19
            assign data_11[m19 + b19*16 + a0*28*16] = data_11_array[a0][b19][m19];
        end
    endgenerate
    generate 
        localparam integer b20 = 20;
        for (m20 = 0; m20 < 16; m20 = m20 + 1) 
        begin: inbit20
            assign data_11[m20 + b20*16 + a0*28*16] = data_11_array[a0][b20][m20];
        end
    endgenerate
    generate 
        localparam integer b21 = 21;
        for (m21 = 0; m21 < 16; m21 = m21 + 1) 
        begin: inbit21
            assign data_11[m21 + b21*16 + a0*28*16] = data_11_array[a0][b21][m21];
        end
    endgenerate
    generate 
        localparam integer b22 = 22;
        for (m22 = 0; m22 < 16; m22 = m22 + 1) 
        begin: inbit22
            assign data_11[m22 + b22*16 + a0*28*16] = data_11_array[a0][b22][m22];
        end
    endgenerate
    generate 
        localparam integer b23 = 23;
        for (m23 = 0; m23 < 16; m23 = m23 + 1) 
        begin: inbit23
            assign data_11[m23 + b23*16 + a0*28*16] = data_11_array[a0][b23][m23];
        end
    endgenerate
    generate 
        localparam integer b24 = 24;
        for (m24 = 0; m24 < 16; m24 = m24 + 1) 
        begin: inbit24
            assign data_11[m24 + b24*16 + a0*28*16] = data_11_array[a0][b24][m24];
        end
    endgenerate
    generate 
        localparam integer b25 = 25;
        for (m25 = 0; m25 < 16; m25 = m25 + 1) 
        begin: inbit25
            assign data_11[m25 + b25*16 + a0*28*16] = data_11_array[a0][b25][m25];
        end
    endgenerate
    generate 
        localparam integer b26 = 26;
        for (m26 = 0; m26 < 16; m26 = m26 + 1) 
        begin: inbit26
            assign data_11[m26 + b26*16 + a0*28*16] = data_11_array[a0][b26][m26];
        end
    endgenerate
    generate 
        localparam integer b27 = 27;
        for (m27 = 0; m27 < 16; m27 = m27 + 1) 
        begin: inbit27
            assign data_11[m27 + b27*16 + a0*28*16] = data_11_array[a0][b27][m27];
        end
    endgenerate
    localparam integer a1 = 1;
    generate 
        localparam integer b28 = 0;
        for (m28 = 0; m28 < 16; m28 = m28 + 1) 
        begin: inbit28
            assign data_11[m28 + b28*16 + a1*28*16] = data_11_array[a1][b28][m28];
        end
    endgenerate
    generate 
        localparam integer b29 = 1;
        for (m29 = 0; m29 < 16; m29 = m29 + 1) 
        begin: inbit29
            assign data_11[m29 + b29*16 + a1*28*16] = data_11_array[a1][b29][m29];
        end
    endgenerate
    generate 
        localparam integer b30 = 2;
        for (m30 = 0; m30 < 16; m30 = m30 + 1) 
        begin: inbit30
            assign data_11[m30 + b30*16 + a1*28*16] = data_11_array[a1][b30][m30];
        end
    endgenerate
    generate 
        localparam integer b31 = 3;
        for (m31 = 0; m31 < 16; m31 = m31 + 1) 
        begin: inbit31
            assign data_11[m31 + b31*16 + a1*28*16] = data_11_array[a1][b31][m31];
        end
    endgenerate
    generate 
        localparam integer b32 = 4;
        for (m32 = 0; m32 < 16; m32 = m32 + 1) 
        begin: inbit32
            assign data_11[m32 + b32*16 + a1*28*16] = data_11_array[a1][b32][m32];
        end
    endgenerate
    generate 
        localparam integer b33 = 5;
        for (m33 = 0; m33 < 16; m33 = m33 + 1) 
        begin: inbit33
            assign data_11[m33 + b33*16 + a1*28*16] = data_11_array[a1][b33][m33];
        end
    endgenerate
    generate 
        localparam integer b34 = 6;
        for (m34 = 0; m34 < 16; m34 = m34 + 1) 
        begin: inbit34
            assign data_11[m34 + b34*16 + a1*28*16] = data_11_array[a1][b34][m34];
        end
    endgenerate
    generate 
        localparam integer b35 = 7;
        for (m35 = 0; m35 < 16; m35 = m35 + 1) 
        begin: inbit35
            assign data_11[m35 + b35*16 + a1*28*16] = data_11_array[a1][b35][m35];
        end
    endgenerate
    generate 
        localparam integer b36 = 8;
        for (m36 = 0; m36 < 16; m36 = m36 + 1) 
        begin: inbit36
            assign data_11[m36 + b36*16 + a1*28*16] = data_11_array[a1][b36][m36];
        end
    endgenerate
    generate 
        localparam integer b37 = 9;
        for (m37 = 0; m37 < 16; m37 = m37 + 1) 
        begin: inbit37
            assign data_11[m37 + b37*16 + a1*28*16] = data_11_array[a1][b37][m37];
        end
    endgenerate
    generate 
        localparam integer b38 = 10;
        for (m38 = 0; m38 < 16; m38 = m38 + 1) 
        begin: inbit38
            assign data_11[m38 + b38*16 + a1*28*16] = data_11_array[a1][b38][m38];
        end
    endgenerate
    generate 
        localparam integer b39 = 11;
        for (m39 = 0; m39 < 16; m39 = m39 + 1) 
        begin: inbit39
            assign data_11[m39 + b39*16 + a1*28*16] = data_11_array[a1][b39][m39];
        end
    endgenerate
    generate 
        localparam integer b40 = 12;
        for (m40 = 0; m40 < 16; m40 = m40 + 1) 
        begin: inbit40
            assign data_11[m40 + b40*16 + a1*28*16] = data_11_array[a1][b40][m40];
        end
    endgenerate
    generate 
        localparam integer b41 = 13;
        for (m41 = 0; m41 < 16; m41 = m41 + 1) 
        begin: inbit41
            assign data_11[m41 + b41*16 + a1*28*16] = data_11_array[a1][b41][m41];
        end
    endgenerate
    generate 
        localparam integer b42 = 14;
        for (m42 = 0; m42 < 16; m42 = m42 + 1) 
        begin: inbit42
            assign data_11[m42 + b42*16 + a1*28*16] = data_11_array[a1][b42][m42];
        end
    endgenerate
    generate 
        localparam integer b43 = 15;
        for (m43 = 0; m43 < 16; m43 = m43 + 1) 
        begin: inbit43
            assign data_11[m43 + b43*16 + a1*28*16] = data_11_array[a1][b43][m43];
        end
    endgenerate
    generate 
        localparam integer b44 = 16;
        for (m44 = 0; m44 < 16; m44 = m44 + 1) 
        begin: inbit44
            assign data_11[m44 + b44*16 + a1*28*16] = data_11_array[a1][b44][m44];
        end
    endgenerate
    generate 
        localparam integer b45 = 17;
        for (m45 = 0; m45 < 16; m45 = m45 + 1) 
        begin: inbit45
            assign data_11[m45 + b45*16 + a1*28*16] = data_11_array[a1][b45][m45];
        end
    endgenerate
    generate 
        localparam integer b46 = 18;
        for (m46 = 0; m46 < 16; m46 = m46 + 1) 
        begin: inbit46
            assign data_11[m46 + b46*16 + a1*28*16] = data_11_array[a1][b46][m46];
        end
    endgenerate
    generate 
        localparam integer b47 = 19;
        for (m47 = 0; m47 < 16; m47 = m47 + 1) 
        begin: inbit47
            assign data_11[m47 + b47*16 + a1*28*16] = data_11_array[a1][b47][m47];
        end
    endgenerate
    generate 
        localparam integer b48 = 20;
        for (m48 = 0; m48 < 16; m48 = m48 + 1) 
        begin: inbit48
            assign data_11[m48 + b48*16 + a1*28*16] = data_11_array[a1][b48][m48];
        end
    endgenerate
    generate 
        localparam integer b49 = 21;
        for (m49 = 0; m49 < 16; m49 = m49 + 1) 
        begin: inbit49
            assign data_11[m49 + b49*16 + a1*28*16] = data_11_array[a1][b49][m49];
        end
    endgenerate
    generate 
        localparam integer b50 = 22;
        for (m50 = 0; m50 < 16; m50 = m50 + 1) 
        begin: inbit50
            assign data_11[m50 + b50*16 + a1*28*16] = data_11_array[a1][b50][m50];
        end
    endgenerate
    generate 
        localparam integer b51 = 23;
        for (m51 = 0; m51 < 16; m51 = m51 + 1) 
        begin: inbit51
            assign data_11[m51 + b51*16 + a1*28*16] = data_11_array[a1][b51][m51];
        end
    endgenerate
    generate 
        localparam integer b52 = 24;
        for (m52 = 0; m52 < 16; m52 = m52 + 1) 
        begin: inbit52
            assign data_11[m52 + b52*16 + a1*28*16] = data_11_array[a1][b52][m52];
        end
    endgenerate
    generate 
        localparam integer b53 = 25;
        for (m53 = 0; m53 < 16; m53 = m53 + 1) 
        begin: inbit53
            assign data_11[m53 + b53*16 + a1*28*16] = data_11_array[a1][b53][m53];
        end
    endgenerate
    generate 
        localparam integer b54 = 26;
        for (m54 = 0; m54 < 16; m54 = m54 + 1) 
        begin: inbit54
            assign data_11[m54 + b54*16 + a1*28*16] = data_11_array[a1][b54][m54];
        end
    endgenerate
    generate 
        localparam integer b55 = 27;
        for (m55 = 0; m55 < 16; m55 = m55 + 1) 
        begin: inbit55
            assign data_11[m55 + b55*16 + a1*28*16] = data_11_array[a1][b55][m55];
        end
    endgenerate
    localparam integer a2 = 2;
    generate 
        localparam integer b56 = 0;
        for (m56 = 0; m56 < 16; m56 = m56 + 1) 
        begin: inbit56
            assign data_11[m56 + b56*16 + a2*28*16] = data_11_array[a2][b56][m56];
        end
    endgenerate
    generate 
        localparam integer b57 = 1;
        for (m57 = 0; m57 < 16; m57 = m57 + 1) 
        begin: inbit57
            assign data_11[m57 + b57*16 + a2*28*16] = data_11_array[a2][b57][m57];
        end
    endgenerate
    generate 
        localparam integer b58 = 2;
        for (m58 = 0; m58 < 16; m58 = m58 + 1) 
        begin: inbit58
            assign data_11[m58 + b58*16 + a2*28*16] = data_11_array[a2][b58][m58];
        end
    endgenerate
    generate 
        localparam integer b59 = 3;
        for (m59 = 0; m59 < 16; m59 = m59 + 1) 
        begin: inbit59
            assign data_11[m59 + b59*16 + a2*28*16] = data_11_array[a2][b59][m59];
        end
    endgenerate
    generate 
        localparam integer b60 = 4;
        for (m60 = 0; m60 < 16; m60 = m60 + 1) 
        begin: inbit60
            assign data_11[m60 + b60*16 + a2*28*16] = data_11_array[a2][b60][m60];
        end
    endgenerate
    generate 
        localparam integer b61 = 5;
        for (m61 = 0; m61 < 16; m61 = m61 + 1) 
        begin: inbit61
            assign data_11[m61 + b61*16 + a2*28*16] = data_11_array[a2][b61][m61];
        end
    endgenerate
    generate 
        localparam integer b62 = 6;
        for (m62 = 0; m62 < 16; m62 = m62 + 1) 
        begin: inbit62
            assign data_11[m62 + b62*16 + a2*28*16] = data_11_array[a2][b62][m62];
        end
    endgenerate
    generate 
        localparam integer b63 = 7;
        for (m63 = 0; m63 < 16; m63 = m63 + 1) 
        begin: inbit63
            assign data_11[m63 + b63*16 + a2*28*16] = data_11_array[a2][b63][m63];
        end
    endgenerate
    generate 
        localparam integer b64 = 8;
        for (m64 = 0; m64 < 16; m64 = m64 + 1) 
        begin: inbit64
            assign data_11[m64 + b64*16 + a2*28*16] = data_11_array[a2][b64][m64];
        end
    endgenerate
    generate 
        localparam integer b65 = 9;
        for (m65 = 0; m65 < 16; m65 = m65 + 1) 
        begin: inbit65
            assign data_11[m65 + b65*16 + a2*28*16] = data_11_array[a2][b65][m65];
        end
    endgenerate
    generate 
        localparam integer b66 = 10;
        for (m66 = 0; m66 < 16; m66 = m66 + 1) 
        begin: inbit66
            assign data_11[m66 + b66*16 + a2*28*16] = data_11_array[a2][b66][m66];
        end
    endgenerate
    generate 
        localparam integer b67 = 11;
        for (m67 = 0; m67 < 16; m67 = m67 + 1) 
        begin: inbit67
            assign data_11[m67 + b67*16 + a2*28*16] = data_11_array[a2][b67][m67];
        end
    endgenerate
    generate 
        localparam integer b68 = 12;
        for (m68 = 0; m68 < 16; m68 = m68 + 1) 
        begin: inbit68
            assign data_11[m68 + b68*16 + a2*28*16] = data_11_array[a2][b68][m68];
        end
    endgenerate
    generate 
        localparam integer b69 = 13;
        for (m69 = 0; m69 < 16; m69 = m69 + 1) 
        begin: inbit69
            assign data_11[m69 + b69*16 + a2*28*16] = data_11_array[a2][b69][m69];
        end
    endgenerate
    generate 
        localparam integer b70 = 14;
        for (m70 = 0; m70 < 16; m70 = m70 + 1) 
        begin: inbit70
            assign data_11[m70 + b70*16 + a2*28*16] = data_11_array[a2][b70][m70];
        end
    endgenerate
    generate 
        localparam integer b71 = 15;
        for (m71 = 0; m71 < 16; m71 = m71 + 1) 
        begin: inbit71
            assign data_11[m71 + b71*16 + a2*28*16] = data_11_array[a2][b71][m71];
        end
    endgenerate
    generate 
        localparam integer b72 = 16;
        for (m72 = 0; m72 < 16; m72 = m72 + 1) 
        begin: inbit72
            assign data_11[m72 + b72*16 + a2*28*16] = data_11_array[a2][b72][m72];
        end
    endgenerate
    generate 
        localparam integer b73 = 17;
        for (m73 = 0; m73 < 16; m73 = m73 + 1) 
        begin: inbit73
            assign data_11[m73 + b73*16 + a2*28*16] = data_11_array[a2][b73][m73];
        end
    endgenerate
    generate 
        localparam integer b74 = 18;
        for (m74 = 0; m74 < 16; m74 = m74 + 1) 
        begin: inbit74
            assign data_11[m74 + b74*16 + a2*28*16] = data_11_array[a2][b74][m74];
        end
    endgenerate
    generate 
        localparam integer b75 = 19;
        for (m75 = 0; m75 < 16; m75 = m75 + 1) 
        begin: inbit75
            assign data_11[m75 + b75*16 + a2*28*16] = data_11_array[a2][b75][m75];
        end
    endgenerate
    generate 
        localparam integer b76 = 20;
        for (m76 = 0; m76 < 16; m76 = m76 + 1) 
        begin: inbit76
            assign data_11[m76 + b76*16 + a2*28*16] = data_11_array[a2][b76][m76];
        end
    endgenerate
    generate 
        localparam integer b77 = 21;
        for (m77 = 0; m77 < 16; m77 = m77 + 1) 
        begin: inbit77
            assign data_11[m77 + b77*16 + a2*28*16] = data_11_array[a2][b77][m77];
        end
    endgenerate
    generate 
        localparam integer b78 = 22;
        for (m78 = 0; m78 < 16; m78 = m78 + 1) 
        begin: inbit78
            assign data_11[m78 + b78*16 + a2*28*16] = data_11_array[a2][b78][m78];
        end
    endgenerate
    generate 
        localparam integer b79 = 23;
        for (m79 = 0; m79 < 16; m79 = m79 + 1) 
        begin: inbit79
            assign data_11[m79 + b79*16 + a2*28*16] = data_11_array[a2][b79][m79];
        end
    endgenerate
    generate 
        localparam integer b80 = 24;
        for (m80 = 0; m80 < 16; m80 = m80 + 1) 
        begin: inbit80
            assign data_11[m80 + b80*16 + a2*28*16] = data_11_array[a2][b80][m80];
        end
    endgenerate
    generate 
        localparam integer b81 = 25;
        for (m81 = 0; m81 < 16; m81 = m81 + 1) 
        begin: inbit81
            assign data_11[m81 + b81*16 + a2*28*16] = data_11_array[a2][b81][m81];
        end
    endgenerate
    generate 
        localparam integer b82 = 26;
        for (m82 = 0; m82 < 16; m82 = m82 + 1) 
        begin: inbit82
            assign data_11[m82 + b82*16 + a2*28*16] = data_11_array[a2][b82][m82];
        end
    endgenerate
    generate 
        localparam integer b83 = 27;
        for (m83 = 0; m83 < 16; m83 = m83 + 1) 
        begin: inbit83
            assign data_11[m83 + b83*16 + a2*28*16] = data_11_array[a2][b83][m83];
        end
    endgenerate
    localparam integer a3 = 3;
    generate 
        localparam integer b84 = 0;
        for (m84 = 0; m84 < 16; m84 = m84 + 1) 
        begin: inbit84
            assign data_11[m84 + b84*16 + a3*28*16] = data_11_array[a3][b84][m84];
        end
    endgenerate
    generate 
        localparam integer b85 = 1;
        for (m85 = 0; m85 < 16; m85 = m85 + 1) 
        begin: inbit85
            assign data_11[m85 + b85*16 + a3*28*16] = data_11_array[a3][b85][m85];
        end
    endgenerate
    generate 
        localparam integer b86 = 2;
        for (m86 = 0; m86 < 16; m86 = m86 + 1) 
        begin: inbit86
            assign data_11[m86 + b86*16 + a3*28*16] = data_11_array[a3][b86][m86];
        end
    endgenerate
    generate 
        localparam integer b87 = 3;
        for (m87 = 0; m87 < 16; m87 = m87 + 1) 
        begin: inbit87
            assign data_11[m87 + b87*16 + a3*28*16] = data_11_array[a3][b87][m87];
        end
    endgenerate
    generate 
        localparam integer b88 = 4;
        for (m88 = 0; m88 < 16; m88 = m88 + 1) 
        begin: inbit88
            assign data_11[m88 + b88*16 + a3*28*16] = data_11_array[a3][b88][m88];
        end
    endgenerate
    generate 
        localparam integer b89 = 5;
        for (m89 = 0; m89 < 16; m89 = m89 + 1) 
        begin: inbit89
            assign data_11[m89 + b89*16 + a3*28*16] = data_11_array[a3][b89][m89];
        end
    endgenerate
    generate 
        localparam integer b90 = 6;
        for (m90 = 0; m90 < 16; m90 = m90 + 1) 
        begin: inbit90
            assign data_11[m90 + b90*16 + a3*28*16] = data_11_array[a3][b90][m90];
        end
    endgenerate
    generate 
        localparam integer b91 = 7;
        for (m91 = 0; m91 < 16; m91 = m91 + 1) 
        begin: inbit91
            assign data_11[m91 + b91*16 + a3*28*16] = data_11_array[a3][b91][m91];
        end
    endgenerate
    generate 
        localparam integer b92 = 8;
        for (m92 = 0; m92 < 16; m92 = m92 + 1) 
        begin: inbit92
            assign data_11[m92 + b92*16 + a3*28*16] = data_11_array[a3][b92][m92];
        end
    endgenerate
    generate 
        localparam integer b93 = 9;
        for (m93 = 0; m93 < 16; m93 = m93 + 1) 
        begin: inbit93
            assign data_11[m93 + b93*16 + a3*28*16] = data_11_array[a3][b93][m93];
        end
    endgenerate
    generate 
        localparam integer b94 = 10;
        for (m94 = 0; m94 < 16; m94 = m94 + 1) 
        begin: inbit94
            assign data_11[m94 + b94*16 + a3*28*16] = data_11_array[a3][b94][m94];
        end
    endgenerate
    generate 
        localparam integer b95 = 11;
        for (m95 = 0; m95 < 16; m95 = m95 + 1) 
        begin: inbit95
            assign data_11[m95 + b95*16 + a3*28*16] = data_11_array[a3][b95][m95];
        end
    endgenerate
    generate 
        localparam integer b96 = 12;
        for (m96 = 0; m96 < 16; m96 = m96 + 1) 
        begin: inbit96
            assign data_11[m96 + b96*16 + a3*28*16] = data_11_array[a3][b96][m96];
        end
    endgenerate
    generate 
        localparam integer b97 = 13;
        for (m97 = 0; m97 < 16; m97 = m97 + 1) 
        begin: inbit97
            assign data_11[m97 + b97*16 + a3*28*16] = data_11_array[a3][b97][m97];
        end
    endgenerate
    generate 
        localparam integer b98 = 14;
        for (m98 = 0; m98 < 16; m98 = m98 + 1) 
        begin: inbit98
            assign data_11[m98 + b98*16 + a3*28*16] = data_11_array[a3][b98][m98];
        end
    endgenerate
    generate 
        localparam integer b99 = 15;
        for (m99 = 0; m99 < 16; m99 = m99 + 1) 
        begin: inbit99
            assign data_11[m99 + b99*16 + a3*28*16] = data_11_array[a3][b99][m99];
        end
    endgenerate
    generate 
        localparam integer b100 = 16;
        for (m100 = 0; m100 < 16; m100 = m100 + 1) 
        begin: inbit100
            assign data_11[m100 + b100*16 + a3*28*16] = data_11_array[a3][b100][m100];
        end
    endgenerate
    generate 
        localparam integer b101 = 17;
        for (m101 = 0; m101 < 16; m101 = m101 + 1) 
        begin: inbit101
            assign data_11[m101 + b101*16 + a3*28*16] = data_11_array[a3][b101][m101];
        end
    endgenerate
    generate 
        localparam integer b102 = 18;
        for (m102 = 0; m102 < 16; m102 = m102 + 1) 
        begin: inbit102
            assign data_11[m102 + b102*16 + a3*28*16] = data_11_array[a3][b102][m102];
        end
    endgenerate
    generate 
        localparam integer b103 = 19;
        for (m103 = 0; m103 < 16; m103 = m103 + 1) 
        begin: inbit103
            assign data_11[m103 + b103*16 + a3*28*16] = data_11_array[a3][b103][m103];
        end
    endgenerate
    generate 
        localparam integer b104 = 20;
        for (m104 = 0; m104 < 16; m104 = m104 + 1) 
        begin: inbit104
            assign data_11[m104 + b104*16 + a3*28*16] = data_11_array[a3][b104][m104];
        end
    endgenerate
    generate 
        localparam integer b105 = 21;
        for (m105 = 0; m105 < 16; m105 = m105 + 1) 
        begin: inbit105
            assign data_11[m105 + b105*16 + a3*28*16] = data_11_array[a3][b105][m105];
        end
    endgenerate
    generate 
        localparam integer b106 = 22;
        for (m106 = 0; m106 < 16; m106 = m106 + 1) 
        begin: inbit106
            assign data_11[m106 + b106*16 + a3*28*16] = data_11_array[a3][b106][m106];
        end
    endgenerate
    generate 
        localparam integer b107 = 23;
        for (m107 = 0; m107 < 16; m107 = m107 + 1) 
        begin: inbit107
            assign data_11[m107 + b107*16 + a3*28*16] = data_11_array[a3][b107][m107];
        end
    endgenerate
    generate 
        localparam integer b108 = 24;
        for (m108 = 0; m108 < 16; m108 = m108 + 1) 
        begin: inbit108
            assign data_11[m108 + b108*16 + a3*28*16] = data_11_array[a3][b108][m108];
        end
    endgenerate
    generate 
        localparam integer b109 = 25;
        for (m109 = 0; m109 < 16; m109 = m109 + 1) 
        begin: inbit109
            assign data_11[m109 + b109*16 + a3*28*16] = data_11_array[a3][b109][m109];
        end
    endgenerate
    generate 
        localparam integer b110 = 26;
        for (m110 = 0; m110 < 16; m110 = m110 + 1) 
        begin: inbit110
            assign data_11[m110 + b110*16 + a3*28*16] = data_11_array[a3][b110][m110];
        end
    endgenerate
    generate 
        localparam integer b111 = 27;
        for (m111 = 0; m111 < 16; m111 = m111 + 1) 
        begin: inbit111
            assign data_11[m111 + b111*16 + a3*28*16] = data_11_array[a3][b111][m111];
        end
    endgenerate
    localparam integer a4 = 4;
    generate 
        localparam integer b112 = 0;
        for (m112 = 0; m112 < 16; m112 = m112 + 1) 
        begin: inbit112
            assign data_11[m112 + b112*16 + a4*28*16] = data_11_array[a4][b112][m112];
        end
    endgenerate
    generate 
        localparam integer b113 = 1;
        for (m113 = 0; m113 < 16; m113 = m113 + 1) 
        begin: inbit113
            assign data_11[m113 + b113*16 + a4*28*16] = data_11_array[a4][b113][m113];
        end
    endgenerate
    generate 
        localparam integer b114 = 2;
        for (m114 = 0; m114 < 16; m114 = m114 + 1) 
        begin: inbit114
            assign data_11[m114 + b114*16 + a4*28*16] = data_11_array[a4][b114][m114];
        end
    endgenerate
    generate 
        localparam integer b115 = 3;
        for (m115 = 0; m115 < 16; m115 = m115 + 1) 
        begin: inbit115
            assign data_11[m115 + b115*16 + a4*28*16] = data_11_array[a4][b115][m115];
        end
    endgenerate
    generate 
        localparam integer b116 = 4;
        for (m116 = 0; m116 < 16; m116 = m116 + 1) 
        begin: inbit116
            assign data_11[m116 + b116*16 + a4*28*16] = data_11_array[a4][b116][m116];
        end
    endgenerate
    generate 
        localparam integer b117 = 5;
        for (m117 = 0; m117 < 16; m117 = m117 + 1) 
        begin: inbit117
            assign data_11[m117 + b117*16 + a4*28*16] = data_11_array[a4][b117][m117];
        end
    endgenerate
    generate 
        localparam integer b118 = 6;
        for (m118 = 0; m118 < 16; m118 = m118 + 1) 
        begin: inbit118
            assign data_11[m118 + b118*16 + a4*28*16] = data_11_array[a4][b118][m118];
        end
    endgenerate
    generate 
        localparam integer b119 = 7;
        for (m119 = 0; m119 < 16; m119 = m119 + 1) 
        begin: inbit119
            assign data_11[m119 + b119*16 + a4*28*16] = data_11_array[a4][b119][m119];
        end
    endgenerate
    generate 
        localparam integer b120 = 8;
        for (m120 = 0; m120 < 16; m120 = m120 + 1) 
        begin: inbit120
            assign data_11[m120 + b120*16 + a4*28*16] = data_11_array[a4][b120][m120];
        end
    endgenerate
    generate 
        localparam integer b121 = 9;
        for (m121 = 0; m121 < 16; m121 = m121 + 1) 
        begin: inbit121
            assign data_11[m121 + b121*16 + a4*28*16] = data_11_array[a4][b121][m121];
        end
    endgenerate
    generate 
        localparam integer b122 = 10;
        for (m122 = 0; m122 < 16; m122 = m122 + 1) 
        begin: inbit122
            assign data_11[m122 + b122*16 + a4*28*16] = data_11_array[a4][b122][m122];
        end
    endgenerate
    generate 
        localparam integer b123 = 11;
        for (m123 = 0; m123 < 16; m123 = m123 + 1) 
        begin: inbit123
            assign data_11[m123 + b123*16 + a4*28*16] = data_11_array[a4][b123][m123];
        end
    endgenerate
    generate 
        localparam integer b124 = 12;
        for (m124 = 0; m124 < 16; m124 = m124 + 1) 
        begin: inbit124
            assign data_11[m124 + b124*16 + a4*28*16] = data_11_array[a4][b124][m124];
        end
    endgenerate
    generate 
        localparam integer b125 = 13;
        for (m125 = 0; m125 < 16; m125 = m125 + 1) 
        begin: inbit125
            assign data_11[m125 + b125*16 + a4*28*16] = data_11_array[a4][b125][m125];
        end
    endgenerate
    generate 
        localparam integer b126 = 14;
        for (m126 = 0; m126 < 16; m126 = m126 + 1) 
        begin: inbit126
            assign data_11[m126 + b126*16 + a4*28*16] = data_11_array[a4][b126][m126];
        end
    endgenerate
    generate 
        localparam integer b127 = 15;
        for (m127 = 0; m127 < 16; m127 = m127 + 1) 
        begin: inbit127
            assign data_11[m127 + b127*16 + a4*28*16] = data_11_array[a4][b127][m127];
        end
    endgenerate
    generate 
        localparam integer b128 = 16;
        for (m128 = 0; m128 < 16; m128 = m128 + 1) 
        begin: inbit128
            assign data_11[m128 + b128*16 + a4*28*16] = data_11_array[a4][b128][m128];
        end
    endgenerate
    generate 
        localparam integer b129 = 17;
        for (m129 = 0; m129 < 16; m129 = m129 + 1) 
        begin: inbit129
            assign data_11[m129 + b129*16 + a4*28*16] = data_11_array[a4][b129][m129];
        end
    endgenerate
    generate 
        localparam integer b130 = 18;
        for (m130 = 0; m130 < 16; m130 = m130 + 1) 
        begin: inbit130
            assign data_11[m130 + b130*16 + a4*28*16] = data_11_array[a4][b130][m130];
        end
    endgenerate
    generate 
        localparam integer b131 = 19;
        for (m131 = 0; m131 < 16; m131 = m131 + 1) 
        begin: inbit131
            assign data_11[m131 + b131*16 + a4*28*16] = data_11_array[a4][b131][m131];
        end
    endgenerate
    generate 
        localparam integer b132 = 20;
        for (m132 = 0; m132 < 16; m132 = m132 + 1) 
        begin: inbit132
            assign data_11[m132 + b132*16 + a4*28*16] = data_11_array[a4][b132][m132];
        end
    endgenerate
    generate 
        localparam integer b133 = 21;
        for (m133 = 0; m133 < 16; m133 = m133 + 1) 
        begin: inbit133
            assign data_11[m133 + b133*16 + a4*28*16] = data_11_array[a4][b133][m133];
        end
    endgenerate
    generate 
        localparam integer b134 = 22;
        for (m134 = 0; m134 < 16; m134 = m134 + 1) 
        begin: inbit134
            assign data_11[m134 + b134*16 + a4*28*16] = data_11_array[a4][b134][m134];
        end
    endgenerate
    generate 
        localparam integer b135 = 23;
        for (m135 = 0; m135 < 16; m135 = m135 + 1) 
        begin: inbit135
            assign data_11[m135 + b135*16 + a4*28*16] = data_11_array[a4][b135][m135];
        end
    endgenerate
    generate 
        localparam integer b136 = 24;
        for (m136 = 0; m136 < 16; m136 = m136 + 1) 
        begin: inbit136
            assign data_11[m136 + b136*16 + a4*28*16] = data_11_array[a4][b136][m136];
        end
    endgenerate
    generate 
        localparam integer b137 = 25;
        for (m137 = 0; m137 < 16; m137 = m137 + 1) 
        begin: inbit137
            assign data_11[m137 + b137*16 + a4*28*16] = data_11_array[a4][b137][m137];
        end
    endgenerate
    generate 
        localparam integer b138 = 26;
        for (m138 = 0; m138 < 16; m138 = m138 + 1) 
        begin: inbit138
            assign data_11[m138 + b138*16 + a4*28*16] = data_11_array[a4][b138][m138];
        end
    endgenerate
    generate 
        localparam integer b139 = 27;
        for (m139 = 0; m139 < 16; m139 = m139 + 1) 
        begin: inbit139
            assign data_11[m139 + b139*16 + a4*28*16] = data_11_array[a4][b139][m139];
        end
    endgenerate
    localparam integer a5 = 5;
    generate 
        localparam integer b140 = 0;
        for (m140 = 0; m140 < 16; m140 = m140 + 1) 
        begin: inbit140
            assign data_11[m140 + b140*16 + a5*28*16] = data_11_array[a5][b140][m140];
        end
    endgenerate
    generate 
        localparam integer b141 = 1;
        for (m141 = 0; m141 < 16; m141 = m141 + 1) 
        begin: inbit141
            assign data_11[m141 + b141*16 + a5*28*16] = data_11_array[a5][b141][m141];
        end
    endgenerate
    generate 
        localparam integer b142 = 2;
        for (m142 = 0; m142 < 16; m142 = m142 + 1) 
        begin: inbit142
            assign data_11[m142 + b142*16 + a5*28*16] = data_11_array[a5][b142][m142];
        end
    endgenerate
    generate 
        localparam integer b143 = 3;
        for (m143 = 0; m143 < 16; m143 = m143 + 1) 
        begin: inbit143
            assign data_11[m143 + b143*16 + a5*28*16] = data_11_array[a5][b143][m143];
        end
    endgenerate
    generate 
        localparam integer b144 = 4;
        for (m144 = 0; m144 < 16; m144 = m144 + 1) 
        begin: inbit144
            assign data_11[m144 + b144*16 + a5*28*16] = data_11_array[a5][b144][m144];
        end
    endgenerate
    generate 
        localparam integer b145 = 5;
        for (m145 = 0; m145 < 16; m145 = m145 + 1) 
        begin: inbit145
            assign data_11[m145 + b145*16 + a5*28*16] = data_11_array[a5][b145][m145];
        end
    endgenerate
    generate 
        localparam integer b146 = 6;
        for (m146 = 0; m146 < 16; m146 = m146 + 1) 
        begin: inbit146
            assign data_11[m146 + b146*16 + a5*28*16] = data_11_array[a5][b146][m146];
        end
    endgenerate
    generate 
        localparam integer b147 = 7;
        for (m147 = 0; m147 < 16; m147 = m147 + 1) 
        begin: inbit147
            assign data_11[m147 + b147*16 + a5*28*16] = data_11_array[a5][b147][m147];
        end
    endgenerate
    generate 
        localparam integer b148 = 8;
        for (m148 = 0; m148 < 16; m148 = m148 + 1) 
        begin: inbit148
            assign data_11[m148 + b148*16 + a5*28*16] = data_11_array[a5][b148][m148];
        end
    endgenerate
    generate 
        localparam integer b149 = 9;
        for (m149 = 0; m149 < 16; m149 = m149 + 1) 
        begin: inbit149
            assign data_11[m149 + b149*16 + a5*28*16] = data_11_array[a5][b149][m149];
        end
    endgenerate
    generate 
        localparam integer b150 = 10;
        for (m150 = 0; m150 < 16; m150 = m150 + 1) 
        begin: inbit150
            assign data_11[m150 + b150*16 + a5*28*16] = data_11_array[a5][b150][m150];
        end
    endgenerate
    generate 
        localparam integer b151 = 11;
        for (m151 = 0; m151 < 16; m151 = m151 + 1) 
        begin: inbit151
            assign data_11[m151 + b151*16 + a5*28*16] = data_11_array[a5][b151][m151];
        end
    endgenerate
    generate 
        localparam integer b152 = 12;
        for (m152 = 0; m152 < 16; m152 = m152 + 1) 
        begin: inbit152
            assign data_11[m152 + b152*16 + a5*28*16] = data_11_array[a5][b152][m152];
        end
    endgenerate
    generate 
        localparam integer b153 = 13;
        for (m153 = 0; m153 < 16; m153 = m153 + 1) 
        begin: inbit153
            assign data_11[m153 + b153*16 + a5*28*16] = data_11_array[a5][b153][m153];
        end
    endgenerate
    generate 
        localparam integer b154 = 14;
        for (m154 = 0; m154 < 16; m154 = m154 + 1) 
        begin: inbit154
            assign data_11[m154 + b154*16 + a5*28*16] = data_11_array[a5][b154][m154];
        end
    endgenerate
    generate 
        localparam integer b155 = 15;
        for (m155 = 0; m155 < 16; m155 = m155 + 1) 
        begin: inbit155
            assign data_11[m155 + b155*16 + a5*28*16] = data_11_array[a5][b155][m155];
        end
    endgenerate
    generate 
        localparam integer b156 = 16;
        for (m156 = 0; m156 < 16; m156 = m156 + 1) 
        begin: inbit156
            assign data_11[m156 + b156*16 + a5*28*16] = data_11_array[a5][b156][m156];
        end
    endgenerate
    generate 
        localparam integer b157 = 17;
        for (m157 = 0; m157 < 16; m157 = m157 + 1) 
        begin: inbit157
            assign data_11[m157 + b157*16 + a5*28*16] = data_11_array[a5][b157][m157];
        end
    endgenerate
    generate 
        localparam integer b158 = 18;
        for (m158 = 0; m158 < 16; m158 = m158 + 1) 
        begin: inbit158
            assign data_11[m158 + b158*16 + a5*28*16] = data_11_array[a5][b158][m158];
        end
    endgenerate
    generate 
        localparam integer b159 = 19;
        for (m159 = 0; m159 < 16; m159 = m159 + 1) 
        begin: inbit159
            assign data_11[m159 + b159*16 + a5*28*16] = data_11_array[a5][b159][m159];
        end
    endgenerate
    generate 
        localparam integer b160 = 20;
        for (m160 = 0; m160 < 16; m160 = m160 + 1) 
        begin: inbit160
            assign data_11[m160 + b160*16 + a5*28*16] = data_11_array[a5][b160][m160];
        end
    endgenerate
    generate 
        localparam integer b161 = 21;
        for (m161 = 0; m161 < 16; m161 = m161 + 1) 
        begin: inbit161
            assign data_11[m161 + b161*16 + a5*28*16] = data_11_array[a5][b161][m161];
        end
    endgenerate
    generate 
        localparam integer b162 = 22;
        for (m162 = 0; m162 < 16; m162 = m162 + 1) 
        begin: inbit162
            assign data_11[m162 + b162*16 + a5*28*16] = data_11_array[a5][b162][m162];
        end
    endgenerate
    generate 
        localparam integer b163 = 23;
        for (m163 = 0; m163 < 16; m163 = m163 + 1) 
        begin: inbit163
            assign data_11[m163 + b163*16 + a5*28*16] = data_11_array[a5][b163][m163];
        end
    endgenerate
    generate 
        localparam integer b164 = 24;
        for (m164 = 0; m164 < 16; m164 = m164 + 1) 
        begin: inbit164
            assign data_11[m164 + b164*16 + a5*28*16] = data_11_array[a5][b164][m164];
        end
    endgenerate
    generate 
        localparam integer b165 = 25;
        for (m165 = 0; m165 < 16; m165 = m165 + 1) 
        begin: inbit165
            assign data_11[m165 + b165*16 + a5*28*16] = data_11_array[a5][b165][m165];
        end
    endgenerate
    generate 
        localparam integer b166 = 26;
        for (m166 = 0; m166 < 16; m166 = m166 + 1) 
        begin: inbit166
            assign data_11[m166 + b166*16 + a5*28*16] = data_11_array[a5][b166][m166];
        end
    endgenerate
    generate 
        localparam integer b167 = 27;
        for (m167 = 0; m167 < 16; m167 = m167 + 1) 
        begin: inbit167
            assign data_11[m167 + b167*16 + a5*28*16] = data_11_array[a5][b167][m167];
        end
    endgenerate
    localparam integer a6 = 6;
    generate 
        localparam integer b168 = 0;
        for (m168 = 0; m168 < 16; m168 = m168 + 1) 
        begin: inbit168
            assign data_11[m168 + b168*16 + a6*28*16] = data_11_array[a6][b168][m168];
        end
    endgenerate
    generate 
        localparam integer b169 = 1;
        for (m169 = 0; m169 < 16; m169 = m169 + 1) 
        begin: inbit169
            assign data_11[m169 + b169*16 + a6*28*16] = data_11_array[a6][b169][m169];
        end
    endgenerate
    generate 
        localparam integer b170 = 2;
        for (m170 = 0; m170 < 16; m170 = m170 + 1) 
        begin: inbit170
            assign data_11[m170 + b170*16 + a6*28*16] = data_11_array[a6][b170][m170];
        end
    endgenerate
    generate 
        localparam integer b171 = 3;
        for (m171 = 0; m171 < 16; m171 = m171 + 1) 
        begin: inbit171
            assign data_11[m171 + b171*16 + a6*28*16] = data_11_array[a6][b171][m171];
        end
    endgenerate
    generate 
        localparam integer b172 = 4;
        for (m172 = 0; m172 < 16; m172 = m172 + 1) 
        begin: inbit172
            assign data_11[m172 + b172*16 + a6*28*16] = data_11_array[a6][b172][m172];
        end
    endgenerate
    generate 
        localparam integer b173 = 5;
        for (m173 = 0; m173 < 16; m173 = m173 + 1) 
        begin: inbit173
            assign data_11[m173 + b173*16 + a6*28*16] = data_11_array[a6][b173][m173];
        end
    endgenerate
    generate 
        localparam integer b174 = 6;
        for (m174 = 0; m174 < 16; m174 = m174 + 1) 
        begin: inbit174
            assign data_11[m174 + b174*16 + a6*28*16] = data_11_array[a6][b174][m174];
        end
    endgenerate
    generate 
        localparam integer b175 = 7;
        for (m175 = 0; m175 < 16; m175 = m175 + 1) 
        begin: inbit175
            assign data_11[m175 + b175*16 + a6*28*16] = data_11_array[a6][b175][m175];
        end
    endgenerate
    generate 
        localparam integer b176 = 8;
        for (m176 = 0; m176 < 16; m176 = m176 + 1) 
        begin: inbit176
            assign data_11[m176 + b176*16 + a6*28*16] = data_11_array[a6][b176][m176];
        end
    endgenerate
    generate 
        localparam integer b177 = 9;
        for (m177 = 0; m177 < 16; m177 = m177 + 1) 
        begin: inbit177
            assign data_11[m177 + b177*16 + a6*28*16] = data_11_array[a6][b177][m177];
        end
    endgenerate
    generate 
        localparam integer b178 = 10;
        for (m178 = 0; m178 < 16; m178 = m178 + 1) 
        begin: inbit178
            assign data_11[m178 + b178*16 + a6*28*16] = data_11_array[a6][b178][m178];
        end
    endgenerate
    generate 
        localparam integer b179 = 11;
        for (m179 = 0; m179 < 16; m179 = m179 + 1) 
        begin: inbit179
            assign data_11[m179 + b179*16 + a6*28*16] = data_11_array[a6][b179][m179];
        end
    endgenerate
    generate 
        localparam integer b180 = 12;
        for (m180 = 0; m180 < 16; m180 = m180 + 1) 
        begin: inbit180
            assign data_11[m180 + b180*16 + a6*28*16] = data_11_array[a6][b180][m180];
        end
    endgenerate
    generate 
        localparam integer b181 = 13;
        for (m181 = 0; m181 < 16; m181 = m181 + 1) 
        begin: inbit181
            assign data_11[m181 + b181*16 + a6*28*16] = data_11_array[a6][b181][m181];
        end
    endgenerate
    generate 
        localparam integer b182 = 14;
        for (m182 = 0; m182 < 16; m182 = m182 + 1) 
        begin: inbit182
            assign data_11[m182 + b182*16 + a6*28*16] = data_11_array[a6][b182][m182];
        end
    endgenerate
    generate 
        localparam integer b183 = 15;
        for (m183 = 0; m183 < 16; m183 = m183 + 1) 
        begin: inbit183
            assign data_11[m183 + b183*16 + a6*28*16] = data_11_array[a6][b183][m183];
        end
    endgenerate
    generate 
        localparam integer b184 = 16;
        for (m184 = 0; m184 < 16; m184 = m184 + 1) 
        begin: inbit184
            assign data_11[m184 + b184*16 + a6*28*16] = data_11_array[a6][b184][m184];
        end
    endgenerate
    generate 
        localparam integer b185 = 17;
        for (m185 = 0; m185 < 16; m185 = m185 + 1) 
        begin: inbit185
            assign data_11[m185 + b185*16 + a6*28*16] = data_11_array[a6][b185][m185];
        end
    endgenerate
    generate 
        localparam integer b186 = 18;
        for (m186 = 0; m186 < 16; m186 = m186 + 1) 
        begin: inbit186
            assign data_11[m186 + b186*16 + a6*28*16] = data_11_array[a6][b186][m186];
        end
    endgenerate
    generate 
        localparam integer b187 = 19;
        for (m187 = 0; m187 < 16; m187 = m187 + 1) 
        begin: inbit187
            assign data_11[m187 + b187*16 + a6*28*16] = data_11_array[a6][b187][m187];
        end
    endgenerate
    generate 
        localparam integer b188 = 20;
        for (m188 = 0; m188 < 16; m188 = m188 + 1) 
        begin: inbit188
            assign data_11[m188 + b188*16 + a6*28*16] = data_11_array[a6][b188][m188];
        end
    endgenerate
    generate 
        localparam integer b189 = 21;
        for (m189 = 0; m189 < 16; m189 = m189 + 1) 
        begin: inbit189
            assign data_11[m189 + b189*16 + a6*28*16] = data_11_array[a6][b189][m189];
        end
    endgenerate
    generate 
        localparam integer b190 = 22;
        for (m190 = 0; m190 < 16; m190 = m190 + 1) 
        begin: inbit190
            assign data_11[m190 + b190*16 + a6*28*16] = data_11_array[a6][b190][m190];
        end
    endgenerate
    generate 
        localparam integer b191 = 23;
        for (m191 = 0; m191 < 16; m191 = m191 + 1) 
        begin: inbit191
            assign data_11[m191 + b191*16 + a6*28*16] = data_11_array[a6][b191][m191];
        end
    endgenerate
    generate 
        localparam integer b192 = 24;
        for (m192 = 0; m192 < 16; m192 = m192 + 1) 
        begin: inbit192
            assign data_11[m192 + b192*16 + a6*28*16] = data_11_array[a6][b192][m192];
        end
    endgenerate
    generate 
        localparam integer b193 = 25;
        for (m193 = 0; m193 < 16; m193 = m193 + 1) 
        begin: inbit193
            assign data_11[m193 + b193*16 + a6*28*16] = data_11_array[a6][b193][m193];
        end
    endgenerate
    generate 
        localparam integer b194 = 26;
        for (m194 = 0; m194 < 16; m194 = m194 + 1) 
        begin: inbit194
            assign data_11[m194 + b194*16 + a6*28*16] = data_11_array[a6][b194][m194];
        end
    endgenerate
    generate 
        localparam integer b195 = 27;
        for (m195 = 0; m195 < 16; m195 = m195 + 1) 
        begin: inbit195
            assign data_11[m195 + b195*16 + a6*28*16] = data_11_array[a6][b195][m195];
        end
    endgenerate
    localparam integer a7 = 7;
    generate 
        localparam integer b196 = 0;
        for (m196 = 0; m196 < 16; m196 = m196 + 1) 
        begin: inbit196
            assign data_11[m196 + b196*16 + a7*28*16] = data_11_array[a7][b196][m196];
        end
    endgenerate
    generate 
        localparam integer b197 = 1;
        for (m197 = 0; m197 < 16; m197 = m197 + 1) 
        begin: inbit197
            assign data_11[m197 + b197*16 + a7*28*16] = data_11_array[a7][b197][m197];
        end
    endgenerate
    generate 
        localparam integer b198 = 2;
        for (m198 = 0; m198 < 16; m198 = m198 + 1) 
        begin: inbit198
            assign data_11[m198 + b198*16 + a7*28*16] = data_11_array[a7][b198][m198];
        end
    endgenerate
    generate 
        localparam integer b199 = 3;
        for (m199 = 0; m199 < 16; m199 = m199 + 1) 
        begin: inbit199
            assign data_11[m199 + b199*16 + a7*28*16] = data_11_array[a7][b199][m199];
        end
    endgenerate
    generate 
        localparam integer b200 = 4;
        for (m200 = 0; m200 < 16; m200 = m200 + 1) 
        begin: inbit200
            assign data_11[m200 + b200*16 + a7*28*16] = data_11_array[a7][b200][m200];
        end
    endgenerate
    generate 
        localparam integer b201 = 5;
        for (m201 = 0; m201 < 16; m201 = m201 + 1) 
        begin: inbit201
            assign data_11[m201 + b201*16 + a7*28*16] = data_11_array[a7][b201][m201];
        end
    endgenerate
    generate 
        localparam integer b202 = 6;
        for (m202 = 0; m202 < 16; m202 = m202 + 1) 
        begin: inbit202
            assign data_11[m202 + b202*16 + a7*28*16] = data_11_array[a7][b202][m202];
        end
    endgenerate
    generate 
        localparam integer b203 = 7;
        for (m203 = 0; m203 < 16; m203 = m203 + 1) 
        begin: inbit203
            assign data_11[m203 + b203*16 + a7*28*16] = data_11_array[a7][b203][m203];
        end
    endgenerate
    generate 
        localparam integer b204 = 8;
        for (m204 = 0; m204 < 16; m204 = m204 + 1) 
        begin: inbit204
            assign data_11[m204 + b204*16 + a7*28*16] = data_11_array[a7][b204][m204];
        end
    endgenerate
    generate 
        localparam integer b205 = 9;
        for (m205 = 0; m205 < 16; m205 = m205 + 1) 
        begin: inbit205
            assign data_11[m205 + b205*16 + a7*28*16] = data_11_array[a7][b205][m205];
        end
    endgenerate
    generate 
        localparam integer b206 = 10;
        for (m206 = 0; m206 < 16; m206 = m206 + 1) 
        begin: inbit206
            assign data_11[m206 + b206*16 + a7*28*16] = data_11_array[a7][b206][m206];
        end
    endgenerate
    generate 
        localparam integer b207 = 11;
        for (m207 = 0; m207 < 16; m207 = m207 + 1) 
        begin: inbit207
            assign data_11[m207 + b207*16 + a7*28*16] = data_11_array[a7][b207][m207];
        end
    endgenerate
    generate 
        localparam integer b208 = 12;
        for (m208 = 0; m208 < 16; m208 = m208 + 1) 
        begin: inbit208
            assign data_11[m208 + b208*16 + a7*28*16] = data_11_array[a7][b208][m208];
        end
    endgenerate
    generate 
        localparam integer b209 = 13;
        for (m209 = 0; m209 < 16; m209 = m209 + 1) 
        begin: inbit209
            assign data_11[m209 + b209*16 + a7*28*16] = data_11_array[a7][b209][m209];
        end
    endgenerate
    generate 
        localparam integer b210 = 14;
        for (m210 = 0; m210 < 16; m210 = m210 + 1) 
        begin: inbit210
            assign data_11[m210 + b210*16 + a7*28*16] = data_11_array[a7][b210][m210];
        end
    endgenerate
    generate 
        localparam integer b211 = 15;
        for (m211 = 0; m211 < 16; m211 = m211 + 1) 
        begin: inbit211
            assign data_11[m211 + b211*16 + a7*28*16] = data_11_array[a7][b211][m211];
        end
    endgenerate
    generate 
        localparam integer b212 = 16;
        for (m212 = 0; m212 < 16; m212 = m212 + 1) 
        begin: inbit212
            assign data_11[m212 + b212*16 + a7*28*16] = data_11_array[a7][b212][m212];
        end
    endgenerate
    generate 
        localparam integer b213 = 17;
        for (m213 = 0; m213 < 16; m213 = m213 + 1) 
        begin: inbit213
            assign data_11[m213 + b213*16 + a7*28*16] = data_11_array[a7][b213][m213];
        end
    endgenerate
    generate 
        localparam integer b214 = 18;
        for (m214 = 0; m214 < 16; m214 = m214 + 1) 
        begin: inbit214
            assign data_11[m214 + b214*16 + a7*28*16] = data_11_array[a7][b214][m214];
        end
    endgenerate
    generate 
        localparam integer b215 = 19;
        for (m215 = 0; m215 < 16; m215 = m215 + 1) 
        begin: inbit215
            assign data_11[m215 + b215*16 + a7*28*16] = data_11_array[a7][b215][m215];
        end
    endgenerate
    generate 
        localparam integer b216 = 20;
        for (m216 = 0; m216 < 16; m216 = m216 + 1) 
        begin: inbit216
            assign data_11[m216 + b216*16 + a7*28*16] = data_11_array[a7][b216][m216];
        end
    endgenerate
    generate 
        localparam integer b217 = 21;
        for (m217 = 0; m217 < 16; m217 = m217 + 1) 
        begin: inbit217
            assign data_11[m217 + b217*16 + a7*28*16] = data_11_array[a7][b217][m217];
        end
    endgenerate
    generate 
        localparam integer b218 = 22;
        for (m218 = 0; m218 < 16; m218 = m218 + 1) 
        begin: inbit218
            assign data_11[m218 + b218*16 + a7*28*16] = data_11_array[a7][b218][m218];
        end
    endgenerate
    generate 
        localparam integer b219 = 23;
        for (m219 = 0; m219 < 16; m219 = m219 + 1) 
        begin: inbit219
            assign data_11[m219 + b219*16 + a7*28*16] = data_11_array[a7][b219][m219];
        end
    endgenerate
    generate 
        localparam integer b220 = 24;
        for (m220 = 0; m220 < 16; m220 = m220 + 1) 
        begin: inbit220
            assign data_11[m220 + b220*16 + a7*28*16] = data_11_array[a7][b220][m220];
        end
    endgenerate
    generate 
        localparam integer b221 = 25;
        for (m221 = 0; m221 < 16; m221 = m221 + 1) 
        begin: inbit221
            assign data_11[m221 + b221*16 + a7*28*16] = data_11_array[a7][b221][m221];
        end
    endgenerate
    generate 
        localparam integer b222 = 26;
        for (m222 = 0; m222 < 16; m222 = m222 + 1) 
        begin: inbit222
            assign data_11[m222 + b222*16 + a7*28*16] = data_11_array[a7][b222][m222];
        end
    endgenerate
    generate 
        localparam integer b223 = 27;
        for (m223 = 0; m223 < 16; m223 = m223 + 1) 
        begin: inbit223
            assign data_11[m223 + b223*16 + a7*28*16] = data_11_array[a7][b223][m223];
        end
    endgenerate
    localparam integer a8 = 8;
    generate 
        localparam integer b224 = 0;
        for (m224 = 0; m224 < 16; m224 = m224 + 1) 
        begin: inbit224
            assign data_11[m224 + b224*16 + a8*28*16] = data_11_array[a8][b224][m224];
        end
    endgenerate
    generate 
        localparam integer b225 = 1;
        for (m225 = 0; m225 < 16; m225 = m225 + 1) 
        begin: inbit225
            assign data_11[m225 + b225*16 + a8*28*16] = data_11_array[a8][b225][m225];
        end
    endgenerate
    generate 
        localparam integer b226 = 2;
        for (m226 = 0; m226 < 16; m226 = m226 + 1) 
        begin: inbit226
            assign data_11[m226 + b226*16 + a8*28*16] = data_11_array[a8][b226][m226];
        end
    endgenerate
    generate 
        localparam integer b227 = 3;
        for (m227 = 0; m227 < 16; m227 = m227 + 1) 
        begin: inbit227
            assign data_11[m227 + b227*16 + a8*28*16] = data_11_array[a8][b227][m227];
        end
    endgenerate
    generate 
        localparam integer b228 = 4;
        for (m228 = 0; m228 < 16; m228 = m228 + 1) 
        begin: inbit228
            assign data_11[m228 + b228*16 + a8*28*16] = data_11_array[a8][b228][m228];
        end
    endgenerate
    generate 
        localparam integer b229 = 5;
        for (m229 = 0; m229 < 16; m229 = m229 + 1) 
        begin: inbit229
            assign data_11[m229 + b229*16 + a8*28*16] = data_11_array[a8][b229][m229];
        end
    endgenerate
    generate 
        localparam integer b230 = 6;
        for (m230 = 0; m230 < 16; m230 = m230 + 1) 
        begin: inbit230
            assign data_11[m230 + b230*16 + a8*28*16] = data_11_array[a8][b230][m230];
        end
    endgenerate
    generate 
        localparam integer b231 = 7;
        for (m231 = 0; m231 < 16; m231 = m231 + 1) 
        begin: inbit231
            assign data_11[m231 + b231*16 + a8*28*16] = data_11_array[a8][b231][m231];
        end
    endgenerate
    generate 
        localparam integer b232 = 8;
        for (m232 = 0; m232 < 16; m232 = m232 + 1) 
        begin: inbit232
            assign data_11[m232 + b232*16 + a8*28*16] = data_11_array[a8][b232][m232];
        end
    endgenerate
    generate 
        localparam integer b233 = 9;
        for (m233 = 0; m233 < 16; m233 = m233 + 1) 
        begin: inbit233
            assign data_11[m233 + b233*16 + a8*28*16] = data_11_array[a8][b233][m233];
        end
    endgenerate
    generate 
        localparam integer b234 = 10;
        for (m234 = 0; m234 < 16; m234 = m234 + 1) 
        begin: inbit234
            assign data_11[m234 + b234*16 + a8*28*16] = data_11_array[a8][b234][m234];
        end
    endgenerate
    generate 
        localparam integer b235 = 11;
        for (m235 = 0; m235 < 16; m235 = m235 + 1) 
        begin: inbit235
            assign data_11[m235 + b235*16 + a8*28*16] = data_11_array[a8][b235][m235];
        end
    endgenerate
    generate 
        localparam integer b236 = 12;
        for (m236 = 0; m236 < 16; m236 = m236 + 1) 
        begin: inbit236
            assign data_11[m236 + b236*16 + a8*28*16] = data_11_array[a8][b236][m236];
        end
    endgenerate
    generate 
        localparam integer b237 = 13;
        for (m237 = 0; m237 < 16; m237 = m237 + 1) 
        begin: inbit237
            assign data_11[m237 + b237*16 + a8*28*16] = data_11_array[a8][b237][m237];
        end
    endgenerate
    generate 
        localparam integer b238 = 14;
        for (m238 = 0; m238 < 16; m238 = m238 + 1) 
        begin: inbit238
            assign data_11[m238 + b238*16 + a8*28*16] = data_11_array[a8][b238][m238];
        end
    endgenerate
    generate 
        localparam integer b239 = 15;
        for (m239 = 0; m239 < 16; m239 = m239 + 1) 
        begin: inbit239
            assign data_11[m239 + b239*16 + a8*28*16] = data_11_array[a8][b239][m239];
        end
    endgenerate
    generate 
        localparam integer b240 = 16;
        for (m240 = 0; m240 < 16; m240 = m240 + 1) 
        begin: inbit240
            assign data_11[m240 + b240*16 + a8*28*16] = data_11_array[a8][b240][m240];
        end
    endgenerate
    generate 
        localparam integer b241 = 17;
        for (m241 = 0; m241 < 16; m241 = m241 + 1) 
        begin: inbit241
            assign data_11[m241 + b241*16 + a8*28*16] = data_11_array[a8][b241][m241];
        end
    endgenerate
    generate 
        localparam integer b242 = 18;
        for (m242 = 0; m242 < 16; m242 = m242 + 1) 
        begin: inbit242
            assign data_11[m242 + b242*16 + a8*28*16] = data_11_array[a8][b242][m242];
        end
    endgenerate
    generate 
        localparam integer b243 = 19;
        for (m243 = 0; m243 < 16; m243 = m243 + 1) 
        begin: inbit243
            assign data_11[m243 + b243*16 + a8*28*16] = data_11_array[a8][b243][m243];
        end
    endgenerate
    generate 
        localparam integer b244 = 20;
        for (m244 = 0; m244 < 16; m244 = m244 + 1) 
        begin: inbit244
            assign data_11[m244 + b244*16 + a8*28*16] = data_11_array[a8][b244][m244];
        end
    endgenerate
    generate 
        localparam integer b245 = 21;
        for (m245 = 0; m245 < 16; m245 = m245 + 1) 
        begin: inbit245
            assign data_11[m245 + b245*16 + a8*28*16] = data_11_array[a8][b245][m245];
        end
    endgenerate
    generate 
        localparam integer b246 = 22;
        for (m246 = 0; m246 < 16; m246 = m246 + 1) 
        begin: inbit246
            assign data_11[m246 + b246*16 + a8*28*16] = data_11_array[a8][b246][m246];
        end
    endgenerate
    generate 
        localparam integer b247 = 23;
        for (m247 = 0; m247 < 16; m247 = m247 + 1) 
        begin: inbit247
            assign data_11[m247 + b247*16 + a8*28*16] = data_11_array[a8][b247][m247];
        end
    endgenerate
    generate 
        localparam integer b248 = 24;
        for (m248 = 0; m248 < 16; m248 = m248 + 1) 
        begin: inbit248
            assign data_11[m248 + b248*16 + a8*28*16] = data_11_array[a8][b248][m248];
        end
    endgenerate
    generate 
        localparam integer b249 = 25;
        for (m249 = 0; m249 < 16; m249 = m249 + 1) 
        begin: inbit249
            assign data_11[m249 + b249*16 + a8*28*16] = data_11_array[a8][b249][m249];
        end
    endgenerate
    generate 
        localparam integer b250 = 26;
        for (m250 = 0; m250 < 16; m250 = m250 + 1) 
        begin: inbit250
            assign data_11[m250 + b250*16 + a8*28*16] = data_11_array[a8][b250][m250];
        end
    endgenerate
    generate 
        localparam integer b251 = 27;
        for (m251 = 0; m251 < 16; m251 = m251 + 1) 
        begin: inbit251
            assign data_11[m251 + b251*16 + a8*28*16] = data_11_array[a8][b251][m251];
        end
    endgenerate
    localparam integer a9 = 9;
    generate 
        localparam integer b252 = 0;
        for (m252 = 0; m252 < 16; m252 = m252 + 1) 
        begin: inbit252
            assign data_11[m252 + b252*16 + a9*28*16] = data_11_array[a9][b252][m252];
        end
    endgenerate
    generate 
        localparam integer b253 = 1;
        for (m253 = 0; m253 < 16; m253 = m253 + 1) 
        begin: inbit253
            assign data_11[m253 + b253*16 + a9*28*16] = data_11_array[a9][b253][m253];
        end
    endgenerate
    generate 
        localparam integer b254 = 2;
        for (m254 = 0; m254 < 16; m254 = m254 + 1) 
        begin: inbit254
            assign data_11[m254 + b254*16 + a9*28*16] = data_11_array[a9][b254][m254];
        end
    endgenerate
    generate 
        localparam integer b255 = 3;
        for (m255 = 0; m255 < 16; m255 = m255 + 1) 
        begin: inbit255
            assign data_11[m255 + b255*16 + a9*28*16] = data_11_array[a9][b255][m255];
        end
    endgenerate
    generate 
        localparam integer b256 = 4;
        for (m256 = 0; m256 < 16; m256 = m256 + 1) 
        begin: inbit256
            assign data_11[m256 + b256*16 + a9*28*16] = data_11_array[a9][b256][m256];
        end
    endgenerate
    generate 
        localparam integer b257 = 5;
        for (m257 = 0; m257 < 16; m257 = m257 + 1) 
        begin: inbit257
            assign data_11[m257 + b257*16 + a9*28*16] = data_11_array[a9][b257][m257];
        end
    endgenerate
    generate 
        localparam integer b258 = 6;
        for (m258 = 0; m258 < 16; m258 = m258 + 1) 
        begin: inbit258
            assign data_11[m258 + b258*16 + a9*28*16] = data_11_array[a9][b258][m258];
        end
    endgenerate
    generate 
        localparam integer b259 = 7;
        for (m259 = 0; m259 < 16; m259 = m259 + 1) 
        begin: inbit259
            assign data_11[m259 + b259*16 + a9*28*16] = data_11_array[a9][b259][m259];
        end
    endgenerate
    generate 
        localparam integer b260 = 8;
        for (m260 = 0; m260 < 16; m260 = m260 + 1) 
        begin: inbit260
            assign data_11[m260 + b260*16 + a9*28*16] = data_11_array[a9][b260][m260];
        end
    endgenerate
    generate 
        localparam integer b261 = 9;
        for (m261 = 0; m261 < 16; m261 = m261 + 1) 
        begin: inbit261
            assign data_11[m261 + b261*16 + a9*28*16] = data_11_array[a9][b261][m261];
        end
    endgenerate
    generate 
        localparam integer b262 = 10;
        for (m262 = 0; m262 < 16; m262 = m262 + 1) 
        begin: inbit262
            assign data_11[m262 + b262*16 + a9*28*16] = data_11_array[a9][b262][m262];
        end
    endgenerate
    generate 
        localparam integer b263 = 11;
        for (m263 = 0; m263 < 16; m263 = m263 + 1) 
        begin: inbit263
            assign data_11[m263 + b263*16 + a9*28*16] = data_11_array[a9][b263][m263];
        end
    endgenerate
    generate 
        localparam integer b264 = 12;
        for (m264 = 0; m264 < 16; m264 = m264 + 1) 
        begin: inbit264
            assign data_11[m264 + b264*16 + a9*28*16] = data_11_array[a9][b264][m264];
        end
    endgenerate
    generate 
        localparam integer b265 = 13;
        for (m265 = 0; m265 < 16; m265 = m265 + 1) 
        begin: inbit265
            assign data_11[m265 + b265*16 + a9*28*16] = data_11_array[a9][b265][m265];
        end
    endgenerate
    generate 
        localparam integer b266 = 14;
        for (m266 = 0; m266 < 16; m266 = m266 + 1) 
        begin: inbit266
            assign data_11[m266 + b266*16 + a9*28*16] = data_11_array[a9][b266][m266];
        end
    endgenerate
    generate 
        localparam integer b267 = 15;
        for (m267 = 0; m267 < 16; m267 = m267 + 1) 
        begin: inbit267
            assign data_11[m267 + b267*16 + a9*28*16] = data_11_array[a9][b267][m267];
        end
    endgenerate
    generate 
        localparam integer b268 = 16;
        for (m268 = 0; m268 < 16; m268 = m268 + 1) 
        begin: inbit268
            assign data_11[m268 + b268*16 + a9*28*16] = data_11_array[a9][b268][m268];
        end
    endgenerate
    generate 
        localparam integer b269 = 17;
        for (m269 = 0; m269 < 16; m269 = m269 + 1) 
        begin: inbit269
            assign data_11[m269 + b269*16 + a9*28*16] = data_11_array[a9][b269][m269];
        end
    endgenerate
    generate 
        localparam integer b270 = 18;
        for (m270 = 0; m270 < 16; m270 = m270 + 1) 
        begin: inbit270
            assign data_11[m270 + b270*16 + a9*28*16] = data_11_array[a9][b270][m270];
        end
    endgenerate
    generate 
        localparam integer b271 = 19;
        for (m271 = 0; m271 < 16; m271 = m271 + 1) 
        begin: inbit271
            assign data_11[m271 + b271*16 + a9*28*16] = data_11_array[a9][b271][m271];
        end
    endgenerate
    generate 
        localparam integer b272 = 20;
        for (m272 = 0; m272 < 16; m272 = m272 + 1) 
        begin: inbit272
            assign data_11[m272 + b272*16 + a9*28*16] = data_11_array[a9][b272][m272];
        end
    endgenerate
    generate 
        localparam integer b273 = 21;
        for (m273 = 0; m273 < 16; m273 = m273 + 1) 
        begin: inbit273
            assign data_11[m273 + b273*16 + a9*28*16] = data_11_array[a9][b273][m273];
        end
    endgenerate
    generate 
        localparam integer b274 = 22;
        for (m274 = 0; m274 < 16; m274 = m274 + 1) 
        begin: inbit274
            assign data_11[m274 + b274*16 + a9*28*16] = data_11_array[a9][b274][m274];
        end
    endgenerate
    generate 
        localparam integer b275 = 23;
        for (m275 = 0; m275 < 16; m275 = m275 + 1) 
        begin: inbit275
            assign data_11[m275 + b275*16 + a9*28*16] = data_11_array[a9][b275][m275];
        end
    endgenerate
    generate 
        localparam integer b276 = 24;
        for (m276 = 0; m276 < 16; m276 = m276 + 1) 
        begin: inbit276
            assign data_11[m276 + b276*16 + a9*28*16] = data_11_array[a9][b276][m276];
        end
    endgenerate
    generate 
        localparam integer b277 = 25;
        for (m277 = 0; m277 < 16; m277 = m277 + 1) 
        begin: inbit277
            assign data_11[m277 + b277*16 + a9*28*16] = data_11_array[a9][b277][m277];
        end
    endgenerate
    generate 
        localparam integer b278 = 26;
        for (m278 = 0; m278 < 16; m278 = m278 + 1) 
        begin: inbit278
            assign data_11[m278 + b278*16 + a9*28*16] = data_11_array[a9][b278][m278];
        end
    endgenerate
    generate 
        localparam integer b279 = 27;
        for (m279 = 0; m279 < 16; m279 = m279 + 1) 
        begin: inbit279
            assign data_11[m279 + b279*16 + a9*28*16] = data_11_array[a9][b279][m279];
        end
    endgenerate
    localparam integer a10 = 10;
    generate 
        localparam integer b280 = 0;
        for (m280 = 0; m280 < 16; m280 = m280 + 1) 
        begin: inbit280
            assign data_11[m280 + b280*16 + a10*28*16] = data_11_array[a10][b280][m280];
        end
    endgenerate
    generate 
        localparam integer b281 = 1;
        for (m281 = 0; m281 < 16; m281 = m281 + 1) 
        begin: inbit281
            assign data_11[m281 + b281*16 + a10*28*16] = data_11_array[a10][b281][m281];
        end
    endgenerate
    generate 
        localparam integer b282 = 2;
        for (m282 = 0; m282 < 16; m282 = m282 + 1) 
        begin: inbit282
            assign data_11[m282 + b282*16 + a10*28*16] = data_11_array[a10][b282][m282];
        end
    endgenerate
    generate 
        localparam integer b283 = 3;
        for (m283 = 0; m283 < 16; m283 = m283 + 1) 
        begin: inbit283
            assign data_11[m283 + b283*16 + a10*28*16] = data_11_array[a10][b283][m283];
        end
    endgenerate
    generate 
        localparam integer b284 = 4;
        for (m284 = 0; m284 < 16; m284 = m284 + 1) 
        begin: inbit284
            assign data_11[m284 + b284*16 + a10*28*16] = data_11_array[a10][b284][m284];
        end
    endgenerate
    generate 
        localparam integer b285 = 5;
        for (m285 = 0; m285 < 16; m285 = m285 + 1) 
        begin: inbit285
            assign data_11[m285 + b285*16 + a10*28*16] = data_11_array[a10][b285][m285];
        end
    endgenerate
    generate 
        localparam integer b286 = 6;
        for (m286 = 0; m286 < 16; m286 = m286 + 1) 
        begin: inbit286
            assign data_11[m286 + b286*16 + a10*28*16] = data_11_array[a10][b286][m286];
        end
    endgenerate
    generate 
        localparam integer b287 = 7;
        for (m287 = 0; m287 < 16; m287 = m287 + 1) 
        begin: inbit287
            assign data_11[m287 + b287*16 + a10*28*16] = data_11_array[a10][b287][m287];
        end
    endgenerate
    generate 
        localparam integer b288 = 8;
        for (m288 = 0; m288 < 16; m288 = m288 + 1) 
        begin: inbit288
            assign data_11[m288 + b288*16 + a10*28*16] = data_11_array[a10][b288][m288];
        end
    endgenerate
    generate 
        localparam integer b289 = 9;
        for (m289 = 0; m289 < 16; m289 = m289 + 1) 
        begin: inbit289
            assign data_11[m289 + b289*16 + a10*28*16] = data_11_array[a10][b289][m289];
        end
    endgenerate
    generate 
        localparam integer b290 = 10;
        for (m290 = 0; m290 < 16; m290 = m290 + 1) 
        begin: inbit290
            assign data_11[m290 + b290*16 + a10*28*16] = data_11_array[a10][b290][m290];
        end
    endgenerate
    generate 
        localparam integer b291 = 11;
        for (m291 = 0; m291 < 16; m291 = m291 + 1) 
        begin: inbit291
            assign data_11[m291 + b291*16 + a10*28*16] = data_11_array[a10][b291][m291];
        end
    endgenerate
    generate 
        localparam integer b292 = 12;
        for (m292 = 0; m292 < 16; m292 = m292 + 1) 
        begin: inbit292
            assign data_11[m292 + b292*16 + a10*28*16] = data_11_array[a10][b292][m292];
        end
    endgenerate
    generate 
        localparam integer b293 = 13;
        for (m293 = 0; m293 < 16; m293 = m293 + 1) 
        begin: inbit293
            assign data_11[m293 + b293*16 + a10*28*16] = data_11_array[a10][b293][m293];
        end
    endgenerate
    generate 
        localparam integer b294 = 14;
        for (m294 = 0; m294 < 16; m294 = m294 + 1) 
        begin: inbit294
            assign data_11[m294 + b294*16 + a10*28*16] = data_11_array[a10][b294][m294];
        end
    endgenerate
    generate 
        localparam integer b295 = 15;
        for (m295 = 0; m295 < 16; m295 = m295 + 1) 
        begin: inbit295
            assign data_11[m295 + b295*16 + a10*28*16] = data_11_array[a10][b295][m295];
        end
    endgenerate
    generate 
        localparam integer b296 = 16;
        for (m296 = 0; m296 < 16; m296 = m296 + 1) 
        begin: inbit296
            assign data_11[m296 + b296*16 + a10*28*16] = data_11_array[a10][b296][m296];
        end
    endgenerate
    generate 
        localparam integer b297 = 17;
        for (m297 = 0; m297 < 16; m297 = m297 + 1) 
        begin: inbit297
            assign data_11[m297 + b297*16 + a10*28*16] = data_11_array[a10][b297][m297];
        end
    endgenerate
    generate 
        localparam integer b298 = 18;
        for (m298 = 0; m298 < 16; m298 = m298 + 1) 
        begin: inbit298
            assign data_11[m298 + b298*16 + a10*28*16] = data_11_array[a10][b298][m298];
        end
    endgenerate
    generate 
        localparam integer b299 = 19;
        for (m299 = 0; m299 < 16; m299 = m299 + 1) 
        begin: inbit299
            assign data_11[m299 + b299*16 + a10*28*16] = data_11_array[a10][b299][m299];
        end
    endgenerate
    generate 
        localparam integer b300 = 20;
        for (m300 = 0; m300 < 16; m300 = m300 + 1) 
        begin: inbit300
            assign data_11[m300 + b300*16 + a10*28*16] = data_11_array[a10][b300][m300];
        end
    endgenerate
    generate 
        localparam integer b301 = 21;
        for (m301 = 0; m301 < 16; m301 = m301 + 1) 
        begin: inbit301
            assign data_11[m301 + b301*16 + a10*28*16] = data_11_array[a10][b301][m301];
        end
    endgenerate
    generate 
        localparam integer b302 = 22;
        for (m302 = 0; m302 < 16; m302 = m302 + 1) 
        begin: inbit302
            assign data_11[m302 + b302*16 + a10*28*16] = data_11_array[a10][b302][m302];
        end
    endgenerate
    generate 
        localparam integer b303 = 23;
        for (m303 = 0; m303 < 16; m303 = m303 + 1) 
        begin: inbit303
            assign data_11[m303 + b303*16 + a10*28*16] = data_11_array[a10][b303][m303];
        end
    endgenerate
    generate 
        localparam integer b304 = 24;
        for (m304 = 0; m304 < 16; m304 = m304 + 1) 
        begin: inbit304
            assign data_11[m304 + b304*16 + a10*28*16] = data_11_array[a10][b304][m304];
        end
    endgenerate
    generate 
        localparam integer b305 = 25;
        for (m305 = 0; m305 < 16; m305 = m305 + 1) 
        begin: inbit305
            assign data_11[m305 + b305*16 + a10*28*16] = data_11_array[a10][b305][m305];
        end
    endgenerate
    generate 
        localparam integer b306 = 26;
        for (m306 = 0; m306 < 16; m306 = m306 + 1) 
        begin: inbit306
            assign data_11[m306 + b306*16 + a10*28*16] = data_11_array[a10][b306][m306];
        end
    endgenerate
    generate 
        localparam integer b307 = 27;
        for (m307 = 0; m307 < 16; m307 = m307 + 1) 
        begin: inbit307
            assign data_11[m307 + b307*16 + a10*28*16] = data_11_array[a10][b307][m307];
        end
    endgenerate
    localparam integer a11 = 11;
    generate 
        localparam integer b308 = 0;
        for (m308 = 0; m308 < 16; m308 = m308 + 1) 
        begin: inbit308
            assign data_11[m308 + b308*16 + a11*28*16] = data_11_array[a11][b308][m308];
        end
    endgenerate
    generate 
        localparam integer b309 = 1;
        for (m309 = 0; m309 < 16; m309 = m309 + 1) 
        begin: inbit309
            assign data_11[m309 + b309*16 + a11*28*16] = data_11_array[a11][b309][m309];
        end
    endgenerate
    generate 
        localparam integer b310 = 2;
        for (m310 = 0; m310 < 16; m310 = m310 + 1) 
        begin: inbit310
            assign data_11[m310 + b310*16 + a11*28*16] = data_11_array[a11][b310][m310];
        end
    endgenerate
    generate 
        localparam integer b311 = 3;
        for (m311 = 0; m311 < 16; m311 = m311 + 1) 
        begin: inbit311
            assign data_11[m311 + b311*16 + a11*28*16] = data_11_array[a11][b311][m311];
        end
    endgenerate
    generate 
        localparam integer b312 = 4;
        for (m312 = 0; m312 < 16; m312 = m312 + 1) 
        begin: inbit312
            assign data_11[m312 + b312*16 + a11*28*16] = data_11_array[a11][b312][m312];
        end
    endgenerate
    generate 
        localparam integer b313 = 5;
        for (m313 = 0; m313 < 16; m313 = m313 + 1) 
        begin: inbit313
            assign data_11[m313 + b313*16 + a11*28*16] = data_11_array[a11][b313][m313];
        end
    endgenerate
    generate 
        localparam integer b314 = 6;
        for (m314 = 0; m314 < 16; m314 = m314 + 1) 
        begin: inbit314
            assign data_11[m314 + b314*16 + a11*28*16] = data_11_array[a11][b314][m314];
        end
    endgenerate
    generate 
        localparam integer b315 = 7;
        for (m315 = 0; m315 < 16; m315 = m315 + 1) 
        begin: inbit315
            assign data_11[m315 + b315*16 + a11*28*16] = data_11_array[a11][b315][m315];
        end
    endgenerate
    generate 
        localparam integer b316 = 8;
        for (m316 = 0; m316 < 16; m316 = m316 + 1) 
        begin: inbit316
            assign data_11[m316 + b316*16 + a11*28*16] = data_11_array[a11][b316][m316];
        end
    endgenerate
    generate 
        localparam integer b317 = 9;
        for (m317 = 0; m317 < 16; m317 = m317 + 1) 
        begin: inbit317
            assign data_11[m317 + b317*16 + a11*28*16] = data_11_array[a11][b317][m317];
        end
    endgenerate
    generate 
        localparam integer b318 = 10;
        for (m318 = 0; m318 < 16; m318 = m318 + 1) 
        begin: inbit318
            assign data_11[m318 + b318*16 + a11*28*16] = data_11_array[a11][b318][m318];
        end
    endgenerate
    generate 
        localparam integer b319 = 11;
        for (m319 = 0; m319 < 16; m319 = m319 + 1) 
        begin: inbit319
            assign data_11[m319 + b319*16 + a11*28*16] = data_11_array[a11][b319][m319];
        end
    endgenerate
    generate 
        localparam integer b320 = 12;
        for (m320 = 0; m320 < 16; m320 = m320 + 1) 
        begin: inbit320
            assign data_11[m320 + b320*16 + a11*28*16] = data_11_array[a11][b320][m320];
        end
    endgenerate
    generate 
        localparam integer b321 = 13;
        for (m321 = 0; m321 < 16; m321 = m321 + 1) 
        begin: inbit321
            assign data_11[m321 + b321*16 + a11*28*16] = data_11_array[a11][b321][m321];
        end
    endgenerate
    generate 
        localparam integer b322 = 14;
        for (m322 = 0; m322 < 16; m322 = m322 + 1) 
        begin: inbit322
            assign data_11[m322 + b322*16 + a11*28*16] = data_11_array[a11][b322][m322];
        end
    endgenerate
    generate 
        localparam integer b323 = 15;
        for (m323 = 0; m323 < 16; m323 = m323 + 1) 
        begin: inbit323
            assign data_11[m323 + b323*16 + a11*28*16] = data_11_array[a11][b323][m323];
        end
    endgenerate
    generate 
        localparam integer b324 = 16;
        for (m324 = 0; m324 < 16; m324 = m324 + 1) 
        begin: inbit324
            assign data_11[m324 + b324*16 + a11*28*16] = data_11_array[a11][b324][m324];
        end
    endgenerate
    generate 
        localparam integer b325 = 17;
        for (m325 = 0; m325 < 16; m325 = m325 + 1) 
        begin: inbit325
            assign data_11[m325 + b325*16 + a11*28*16] = data_11_array[a11][b325][m325];
        end
    endgenerate
    generate 
        localparam integer b326 = 18;
        for (m326 = 0; m326 < 16; m326 = m326 + 1) 
        begin: inbit326
            assign data_11[m326 + b326*16 + a11*28*16] = data_11_array[a11][b326][m326];
        end
    endgenerate
    generate 
        localparam integer b327 = 19;
        for (m327 = 0; m327 < 16; m327 = m327 + 1) 
        begin: inbit327
            assign data_11[m327 + b327*16 + a11*28*16] = data_11_array[a11][b327][m327];
        end
    endgenerate
    generate 
        localparam integer b328 = 20;
        for (m328 = 0; m328 < 16; m328 = m328 + 1) 
        begin: inbit328
            assign data_11[m328 + b328*16 + a11*28*16] = data_11_array[a11][b328][m328];
        end
    endgenerate
    generate 
        localparam integer b329 = 21;
        for (m329 = 0; m329 < 16; m329 = m329 + 1) 
        begin: inbit329
            assign data_11[m329 + b329*16 + a11*28*16] = data_11_array[a11][b329][m329];
        end
    endgenerate
    generate 
        localparam integer b330 = 22;
        for (m330 = 0; m330 < 16; m330 = m330 + 1) 
        begin: inbit330
            assign data_11[m330 + b330*16 + a11*28*16] = data_11_array[a11][b330][m330];
        end
    endgenerate
    generate 
        localparam integer b331 = 23;
        for (m331 = 0; m331 < 16; m331 = m331 + 1) 
        begin: inbit331
            assign data_11[m331 + b331*16 + a11*28*16] = data_11_array[a11][b331][m331];
        end
    endgenerate
    generate 
        localparam integer b332 = 24;
        for (m332 = 0; m332 < 16; m332 = m332 + 1) 
        begin: inbit332
            assign data_11[m332 + b332*16 + a11*28*16] = data_11_array[a11][b332][m332];
        end
    endgenerate
    generate 
        localparam integer b333 = 25;
        for (m333 = 0; m333 < 16; m333 = m333 + 1) 
        begin: inbit333
            assign data_11[m333 + b333*16 + a11*28*16] = data_11_array[a11][b333][m333];
        end
    endgenerate
    generate 
        localparam integer b334 = 26;
        for (m334 = 0; m334 < 16; m334 = m334 + 1) 
        begin: inbit334
            assign data_11[m334 + b334*16 + a11*28*16] = data_11_array[a11][b334][m334];
        end
    endgenerate
    generate 
        localparam integer b335 = 27;
        for (m335 = 0; m335 < 16; m335 = m335 + 1) 
        begin: inbit335
            assign data_11[m335 + b335*16 + a11*28*16] = data_11_array[a11][b335][m335];
        end
    endgenerate
    localparam integer a12 = 12;
    generate 
        localparam integer b336 = 0;
        for (m336 = 0; m336 < 16; m336 = m336 + 1) 
        begin: inbit336
            assign data_11[m336 + b336*16 + a12*28*16] = data_11_array[a12][b336][m336];
        end
    endgenerate
    generate 
        localparam integer b337 = 1;
        for (m337 = 0; m337 < 16; m337 = m337 + 1) 
        begin: inbit337
            assign data_11[m337 + b337*16 + a12*28*16] = data_11_array[a12][b337][m337];
        end
    endgenerate
    generate 
        localparam integer b338 = 2;
        for (m338 = 0; m338 < 16; m338 = m338 + 1) 
        begin: inbit338
            assign data_11[m338 + b338*16 + a12*28*16] = data_11_array[a12][b338][m338];
        end
    endgenerate
    generate 
        localparam integer b339 = 3;
        for (m339 = 0; m339 < 16; m339 = m339 + 1) 
        begin: inbit339
            assign data_11[m339 + b339*16 + a12*28*16] = data_11_array[a12][b339][m339];
        end
    endgenerate
    generate 
        localparam integer b340 = 4;
        for (m340 = 0; m340 < 16; m340 = m340 + 1) 
        begin: inbit340
            assign data_11[m340 + b340*16 + a12*28*16] = data_11_array[a12][b340][m340];
        end
    endgenerate
    generate 
        localparam integer b341 = 5;
        for (m341 = 0; m341 < 16; m341 = m341 + 1) 
        begin: inbit341
            assign data_11[m341 + b341*16 + a12*28*16] = data_11_array[a12][b341][m341];
        end
    endgenerate
    generate 
        localparam integer b342 = 6;
        for (m342 = 0; m342 < 16; m342 = m342 + 1) 
        begin: inbit342
            assign data_11[m342 + b342*16 + a12*28*16] = data_11_array[a12][b342][m342];
        end
    endgenerate
    generate 
        localparam integer b343 = 7;
        for (m343 = 0; m343 < 16; m343 = m343 + 1) 
        begin: inbit343
            assign data_11[m343 + b343*16 + a12*28*16] = data_11_array[a12][b343][m343];
        end
    endgenerate
    generate 
        localparam integer b344 = 8;
        for (m344 = 0; m344 < 16; m344 = m344 + 1) 
        begin: inbit344
            assign data_11[m344 + b344*16 + a12*28*16] = data_11_array[a12][b344][m344];
        end
    endgenerate
    generate 
        localparam integer b345 = 9;
        for (m345 = 0; m345 < 16; m345 = m345 + 1) 
        begin: inbit345
            assign data_11[m345 + b345*16 + a12*28*16] = data_11_array[a12][b345][m345];
        end
    endgenerate
    generate 
        localparam integer b346 = 10;
        for (m346 = 0; m346 < 16; m346 = m346 + 1) 
        begin: inbit346
            assign data_11[m346 + b346*16 + a12*28*16] = data_11_array[a12][b346][m346];
        end
    endgenerate
    generate 
        localparam integer b347 = 11;
        for (m347 = 0; m347 < 16; m347 = m347 + 1) 
        begin: inbit347
            assign data_11[m347 + b347*16 + a12*28*16] = data_11_array[a12][b347][m347];
        end
    endgenerate
    generate 
        localparam integer b348 = 12;
        for (m348 = 0; m348 < 16; m348 = m348 + 1) 
        begin: inbit348
            assign data_11[m348 + b348*16 + a12*28*16] = data_11_array[a12][b348][m348];
        end
    endgenerate
    generate 
        localparam integer b349 = 13;
        for (m349 = 0; m349 < 16; m349 = m349 + 1) 
        begin: inbit349
            assign data_11[m349 + b349*16 + a12*28*16] = data_11_array[a12][b349][m349];
        end
    endgenerate
    generate 
        localparam integer b350 = 14;
        for (m350 = 0; m350 < 16; m350 = m350 + 1) 
        begin: inbit350
            assign data_11[m350 + b350*16 + a12*28*16] = data_11_array[a12][b350][m350];
        end
    endgenerate
    generate 
        localparam integer b351 = 15;
        for (m351 = 0; m351 < 16; m351 = m351 + 1) 
        begin: inbit351
            assign data_11[m351 + b351*16 + a12*28*16] = data_11_array[a12][b351][m351];
        end
    endgenerate
    generate 
        localparam integer b352 = 16;
        for (m352 = 0; m352 < 16; m352 = m352 + 1) 
        begin: inbit352
            assign data_11[m352 + b352*16 + a12*28*16] = data_11_array[a12][b352][m352];
        end
    endgenerate
    generate 
        localparam integer b353 = 17;
        for (m353 = 0; m353 < 16; m353 = m353 + 1) 
        begin: inbit353
            assign data_11[m353 + b353*16 + a12*28*16] = data_11_array[a12][b353][m353];
        end
    endgenerate
    generate 
        localparam integer b354 = 18;
        for (m354 = 0; m354 < 16; m354 = m354 + 1) 
        begin: inbit354
            assign data_11[m354 + b354*16 + a12*28*16] = data_11_array[a12][b354][m354];
        end
    endgenerate
    generate 
        localparam integer b355 = 19;
        for (m355 = 0; m355 < 16; m355 = m355 + 1) 
        begin: inbit355
            assign data_11[m355 + b355*16 + a12*28*16] = data_11_array[a12][b355][m355];
        end
    endgenerate
    generate 
        localparam integer b356 = 20;
        for (m356 = 0; m356 < 16; m356 = m356 + 1) 
        begin: inbit356
            assign data_11[m356 + b356*16 + a12*28*16] = data_11_array[a12][b356][m356];
        end
    endgenerate
    generate 
        localparam integer b357 = 21;
        for (m357 = 0; m357 < 16; m357 = m357 + 1) 
        begin: inbit357
            assign data_11[m357 + b357*16 + a12*28*16] = data_11_array[a12][b357][m357];
        end
    endgenerate
    generate 
        localparam integer b358 = 22;
        for (m358 = 0; m358 < 16; m358 = m358 + 1) 
        begin: inbit358
            assign data_11[m358 + b358*16 + a12*28*16] = data_11_array[a12][b358][m358];
        end
    endgenerate
    generate 
        localparam integer b359 = 23;
        for (m359 = 0; m359 < 16; m359 = m359 + 1) 
        begin: inbit359
            assign data_11[m359 + b359*16 + a12*28*16] = data_11_array[a12][b359][m359];
        end
    endgenerate
    generate 
        localparam integer b360 = 24;
        for (m360 = 0; m360 < 16; m360 = m360 + 1) 
        begin: inbit360
            assign data_11[m360 + b360*16 + a12*28*16] = data_11_array[a12][b360][m360];
        end
    endgenerate
    generate 
        localparam integer b361 = 25;
        for (m361 = 0; m361 < 16; m361 = m361 + 1) 
        begin: inbit361
            assign data_11[m361 + b361*16 + a12*28*16] = data_11_array[a12][b361][m361];
        end
    endgenerate
    generate 
        localparam integer b362 = 26;
        for (m362 = 0; m362 < 16; m362 = m362 + 1) 
        begin: inbit362
            assign data_11[m362 + b362*16 + a12*28*16] = data_11_array[a12][b362][m362];
        end
    endgenerate
    generate 
        localparam integer b363 = 27;
        for (m363 = 0; m363 < 16; m363 = m363 + 1) 
        begin: inbit363
            assign data_11[m363 + b363*16 + a12*28*16] = data_11_array[a12][b363][m363];
        end
    endgenerate
    localparam integer a13 = 13;
    generate 
        localparam integer b364 = 0;
        for (m364 = 0; m364 < 16; m364 = m364 + 1) 
        begin: inbit364
            assign data_11[m364 + b364*16 + a13*28*16] = data_11_array[a13][b364][m364];
        end
    endgenerate
    generate 
        localparam integer b365 = 1;
        for (m365 = 0; m365 < 16; m365 = m365 + 1) 
        begin: inbit365
            assign data_11[m365 + b365*16 + a13*28*16] = data_11_array[a13][b365][m365];
        end
    endgenerate
    generate 
        localparam integer b366 = 2;
        for (m366 = 0; m366 < 16; m366 = m366 + 1) 
        begin: inbit366
            assign data_11[m366 + b366*16 + a13*28*16] = data_11_array[a13][b366][m366];
        end
    endgenerate
    generate 
        localparam integer b367 = 3;
        for (m367 = 0; m367 < 16; m367 = m367 + 1) 
        begin: inbit367
            assign data_11[m367 + b367*16 + a13*28*16] = data_11_array[a13][b367][m367];
        end
    endgenerate
    generate 
        localparam integer b368 = 4;
        for (m368 = 0; m368 < 16; m368 = m368 + 1) 
        begin: inbit368
            assign data_11[m368 + b368*16 + a13*28*16] = data_11_array[a13][b368][m368];
        end
    endgenerate
    generate 
        localparam integer b369 = 5;
        for (m369 = 0; m369 < 16; m369 = m369 + 1) 
        begin: inbit369
            assign data_11[m369 + b369*16 + a13*28*16] = data_11_array[a13][b369][m369];
        end
    endgenerate
    generate 
        localparam integer b370 = 6;
        for (m370 = 0; m370 < 16; m370 = m370 + 1) 
        begin: inbit370
            assign data_11[m370 + b370*16 + a13*28*16] = data_11_array[a13][b370][m370];
        end
    endgenerate
    generate 
        localparam integer b371 = 7;
        for (m371 = 0; m371 < 16; m371 = m371 + 1) 
        begin: inbit371
            assign data_11[m371 + b371*16 + a13*28*16] = data_11_array[a13][b371][m371];
        end
    endgenerate
    generate 
        localparam integer b372 = 8;
        for (m372 = 0; m372 < 16; m372 = m372 + 1) 
        begin: inbit372
            assign data_11[m372 + b372*16 + a13*28*16] = data_11_array[a13][b372][m372];
        end
    endgenerate
    generate 
        localparam integer b373 = 9;
        for (m373 = 0; m373 < 16; m373 = m373 + 1) 
        begin: inbit373
            assign data_11[m373 + b373*16 + a13*28*16] = data_11_array[a13][b373][m373];
        end
    endgenerate
    generate 
        localparam integer b374 = 10;
        for (m374 = 0; m374 < 16; m374 = m374 + 1) 
        begin: inbit374
            assign data_11[m374 + b374*16 + a13*28*16] = data_11_array[a13][b374][m374];
        end
    endgenerate
    generate 
        localparam integer b375 = 11;
        for (m375 = 0; m375 < 16; m375 = m375 + 1) 
        begin: inbit375
            assign data_11[m375 + b375*16 + a13*28*16] = data_11_array[a13][b375][m375];
        end
    endgenerate
    generate 
        localparam integer b376 = 12;
        for (m376 = 0; m376 < 16; m376 = m376 + 1) 
        begin: inbit376
            assign data_11[m376 + b376*16 + a13*28*16] = data_11_array[a13][b376][m376];
        end
    endgenerate
    generate 
        localparam integer b377 = 13;
        for (m377 = 0; m377 < 16; m377 = m377 + 1) 
        begin: inbit377
            assign data_11[m377 + b377*16 + a13*28*16] = data_11_array[a13][b377][m377];
        end
    endgenerate
    generate 
        localparam integer b378 = 14;
        for (m378 = 0; m378 < 16; m378 = m378 + 1) 
        begin: inbit378
            assign data_11[m378 + b378*16 + a13*28*16] = data_11_array[a13][b378][m378];
        end
    endgenerate
    generate 
        localparam integer b379 = 15;
        for (m379 = 0; m379 < 16; m379 = m379 + 1) 
        begin: inbit379
            assign data_11[m379 + b379*16 + a13*28*16] = data_11_array[a13][b379][m379];
        end
    endgenerate
    generate 
        localparam integer b380 = 16;
        for (m380 = 0; m380 < 16; m380 = m380 + 1) 
        begin: inbit380
            assign data_11[m380 + b380*16 + a13*28*16] = data_11_array[a13][b380][m380];
        end
    endgenerate
    generate 
        localparam integer b381 = 17;
        for (m381 = 0; m381 < 16; m381 = m381 + 1) 
        begin: inbit381
            assign data_11[m381 + b381*16 + a13*28*16] = data_11_array[a13][b381][m381];
        end
    endgenerate
    generate 
        localparam integer b382 = 18;
        for (m382 = 0; m382 < 16; m382 = m382 + 1) 
        begin: inbit382
            assign data_11[m382 + b382*16 + a13*28*16] = data_11_array[a13][b382][m382];
        end
    endgenerate
    generate 
        localparam integer b383 = 19;
        for (m383 = 0; m383 < 16; m383 = m383 + 1) 
        begin: inbit383
            assign data_11[m383 + b383*16 + a13*28*16] = data_11_array[a13][b383][m383];
        end
    endgenerate
    generate 
        localparam integer b384 = 20;
        for (m384 = 0; m384 < 16; m384 = m384 + 1) 
        begin: inbit384
            assign data_11[m384 + b384*16 + a13*28*16] = data_11_array[a13][b384][m384];
        end
    endgenerate
    generate 
        localparam integer b385 = 21;
        for (m385 = 0; m385 < 16; m385 = m385 + 1) 
        begin: inbit385
            assign data_11[m385 + b385*16 + a13*28*16] = data_11_array[a13][b385][m385];
        end
    endgenerate
    generate 
        localparam integer b386 = 22;
        for (m386 = 0; m386 < 16; m386 = m386 + 1) 
        begin: inbit386
            assign data_11[m386 + b386*16 + a13*28*16] = data_11_array[a13][b386][m386];
        end
    endgenerate
    generate 
        localparam integer b387 = 23;
        for (m387 = 0; m387 < 16; m387 = m387 + 1) 
        begin: inbit387
            assign data_11[m387 + b387*16 + a13*28*16] = data_11_array[a13][b387][m387];
        end
    endgenerate
    generate 
        localparam integer b388 = 24;
        for (m388 = 0; m388 < 16; m388 = m388 + 1) 
        begin: inbit388
            assign data_11[m388 + b388*16 + a13*28*16] = data_11_array[a13][b388][m388];
        end
    endgenerate
    generate 
        localparam integer b389 = 25;
        for (m389 = 0; m389 < 16; m389 = m389 + 1) 
        begin: inbit389
            assign data_11[m389 + b389*16 + a13*28*16] = data_11_array[a13][b389][m389];
        end
    endgenerate
    generate 
        localparam integer b390 = 26;
        for (m390 = 0; m390 < 16; m390 = m390 + 1) 
        begin: inbit390
            assign data_11[m390 + b390*16 + a13*28*16] = data_11_array[a13][b390][m390];
        end
    endgenerate
    generate 
        localparam integer b391 = 27;
        for (m391 = 0; m391 < 16; m391 = m391 + 1) 
        begin: inbit391
            assign data_11[m391 + b391*16 + a13*28*16] = data_11_array[a13][b391][m391];
        end
    endgenerate
    localparam integer a14 = 14;
    generate 
        localparam integer b392 = 0;
        for (m392 = 0; m392 < 16; m392 = m392 + 1) 
        begin: inbit392
            assign data_11[m392 + b392*16 + a14*28*16] = data_11_array[a14][b392][m392];
        end
    endgenerate
    generate 
        localparam integer b393 = 1;
        for (m393 = 0; m393 < 16; m393 = m393 + 1) 
        begin: inbit393
            assign data_11[m393 + b393*16 + a14*28*16] = data_11_array[a14][b393][m393];
        end
    endgenerate
    generate 
        localparam integer b394 = 2;
        for (m394 = 0; m394 < 16; m394 = m394 + 1) 
        begin: inbit394
            assign data_11[m394 + b394*16 + a14*28*16] = data_11_array[a14][b394][m394];
        end
    endgenerate
    generate 
        localparam integer b395 = 3;
        for (m395 = 0; m395 < 16; m395 = m395 + 1) 
        begin: inbit395
            assign data_11[m395 + b395*16 + a14*28*16] = data_11_array[a14][b395][m395];
        end
    endgenerate
    generate 
        localparam integer b396 = 4;
        for (m396 = 0; m396 < 16; m396 = m396 + 1) 
        begin: inbit396
            assign data_11[m396 + b396*16 + a14*28*16] = data_11_array[a14][b396][m396];
        end
    endgenerate
    generate 
        localparam integer b397 = 5;
        for (m397 = 0; m397 < 16; m397 = m397 + 1) 
        begin: inbit397
            assign data_11[m397 + b397*16 + a14*28*16] = data_11_array[a14][b397][m397];
        end
    endgenerate
    generate 
        localparam integer b398 = 6;
        for (m398 = 0; m398 < 16; m398 = m398 + 1) 
        begin: inbit398
            assign data_11[m398 + b398*16 + a14*28*16] = data_11_array[a14][b398][m398];
        end
    endgenerate
    generate 
        localparam integer b399 = 7;
        for (m399 = 0; m399 < 16; m399 = m399 + 1) 
        begin: inbit399
            assign data_11[m399 + b399*16 + a14*28*16] = data_11_array[a14][b399][m399];
        end
    endgenerate
    generate 
        localparam integer b400 = 8;
        for (m400 = 0; m400 < 16; m400 = m400 + 1) 
        begin: inbit400
            assign data_11[m400 + b400*16 + a14*28*16] = data_11_array[a14][b400][m400];
        end
    endgenerate
    generate 
        localparam integer b401 = 9;
        for (m401 = 0; m401 < 16; m401 = m401 + 1) 
        begin: inbit401
            assign data_11[m401 + b401*16 + a14*28*16] = data_11_array[a14][b401][m401];
        end
    endgenerate
    generate 
        localparam integer b402 = 10;
        for (m402 = 0; m402 < 16; m402 = m402 + 1) 
        begin: inbit402
            assign data_11[m402 + b402*16 + a14*28*16] = data_11_array[a14][b402][m402];
        end
    endgenerate
    generate 
        localparam integer b403 = 11;
        for (m403 = 0; m403 < 16; m403 = m403 + 1) 
        begin: inbit403
            assign data_11[m403 + b403*16 + a14*28*16] = data_11_array[a14][b403][m403];
        end
    endgenerate
    generate 
        localparam integer b404 = 12;
        for (m404 = 0; m404 < 16; m404 = m404 + 1) 
        begin: inbit404
            assign data_11[m404 + b404*16 + a14*28*16] = data_11_array[a14][b404][m404];
        end
    endgenerate
    generate 
        localparam integer b405 = 13;
        for (m405 = 0; m405 < 16; m405 = m405 + 1) 
        begin: inbit405
            assign data_11[m405 + b405*16 + a14*28*16] = data_11_array[a14][b405][m405];
        end
    endgenerate
    generate 
        localparam integer b406 = 14;
        for (m406 = 0; m406 < 16; m406 = m406 + 1) 
        begin: inbit406
            assign data_11[m406 + b406*16 + a14*28*16] = data_11_array[a14][b406][m406];
        end
    endgenerate
    generate 
        localparam integer b407 = 15;
        for (m407 = 0; m407 < 16; m407 = m407 + 1) 
        begin: inbit407
            assign data_11[m407 + b407*16 + a14*28*16] = data_11_array[a14][b407][m407];
        end
    endgenerate
    generate 
        localparam integer b408 = 16;
        for (m408 = 0; m408 < 16; m408 = m408 + 1) 
        begin: inbit408
            assign data_11[m408 + b408*16 + a14*28*16] = data_11_array[a14][b408][m408];
        end
    endgenerate
    generate 
        localparam integer b409 = 17;
        for (m409 = 0; m409 < 16; m409 = m409 + 1) 
        begin: inbit409
            assign data_11[m409 + b409*16 + a14*28*16] = data_11_array[a14][b409][m409];
        end
    endgenerate
    generate 
        localparam integer b410 = 18;
        for (m410 = 0; m410 < 16; m410 = m410 + 1) 
        begin: inbit410
            assign data_11[m410 + b410*16 + a14*28*16] = data_11_array[a14][b410][m410];
        end
    endgenerate
    generate 
        localparam integer b411 = 19;
        for (m411 = 0; m411 < 16; m411 = m411 + 1) 
        begin: inbit411
            assign data_11[m411 + b411*16 + a14*28*16] = data_11_array[a14][b411][m411];
        end
    endgenerate
    generate 
        localparam integer b412 = 20;
        for (m412 = 0; m412 < 16; m412 = m412 + 1) 
        begin: inbit412
            assign data_11[m412 + b412*16 + a14*28*16] = data_11_array[a14][b412][m412];
        end
    endgenerate
    generate 
        localparam integer b413 = 21;
        for (m413 = 0; m413 < 16; m413 = m413 + 1) 
        begin: inbit413
            assign data_11[m413 + b413*16 + a14*28*16] = data_11_array[a14][b413][m413];
        end
    endgenerate
    generate 
        localparam integer b414 = 22;
        for (m414 = 0; m414 < 16; m414 = m414 + 1) 
        begin: inbit414
            assign data_11[m414 + b414*16 + a14*28*16] = data_11_array[a14][b414][m414];
        end
    endgenerate
    generate 
        localparam integer b415 = 23;
        for (m415 = 0; m415 < 16; m415 = m415 + 1) 
        begin: inbit415
            assign data_11[m415 + b415*16 + a14*28*16] = data_11_array[a14][b415][m415];
        end
    endgenerate
    generate 
        localparam integer b416 = 24;
        for (m416 = 0; m416 < 16; m416 = m416 + 1) 
        begin: inbit416
            assign data_11[m416 + b416*16 + a14*28*16] = data_11_array[a14][b416][m416];
        end
    endgenerate
    generate 
        localparam integer b417 = 25;
        for (m417 = 0; m417 < 16; m417 = m417 + 1) 
        begin: inbit417
            assign data_11[m417 + b417*16 + a14*28*16] = data_11_array[a14][b417][m417];
        end
    endgenerate
    generate 
        localparam integer b418 = 26;
        for (m418 = 0; m418 < 16; m418 = m418 + 1) 
        begin: inbit418
            assign data_11[m418 + b418*16 + a14*28*16] = data_11_array[a14][b418][m418];
        end
    endgenerate
    generate 
        localparam integer b419 = 27;
        for (m419 = 0; m419 < 16; m419 = m419 + 1) 
        begin: inbit419
            assign data_11[m419 + b419*16 + a14*28*16] = data_11_array[a14][b419][m419];
        end
    endgenerate
    localparam integer a15 = 15;
    generate 
        localparam integer b420 = 0;
        for (m420 = 0; m420 < 16; m420 = m420 + 1) 
        begin: inbit420
            assign data_11[m420 + b420*16 + a15*28*16] = data_11_array[a15][b420][m420];
        end
    endgenerate
    generate 
        localparam integer b421 = 1;
        for (m421 = 0; m421 < 16; m421 = m421 + 1) 
        begin: inbit421
            assign data_11[m421 + b421*16 + a15*28*16] = data_11_array[a15][b421][m421];
        end
    endgenerate
    generate 
        localparam integer b422 = 2;
        for (m422 = 0; m422 < 16; m422 = m422 + 1) 
        begin: inbit422
            assign data_11[m422 + b422*16 + a15*28*16] = data_11_array[a15][b422][m422];
        end
    endgenerate
    generate 
        localparam integer b423 = 3;
        for (m423 = 0; m423 < 16; m423 = m423 + 1) 
        begin: inbit423
            assign data_11[m423 + b423*16 + a15*28*16] = data_11_array[a15][b423][m423];
        end
    endgenerate
    generate 
        localparam integer b424 = 4;
        for (m424 = 0; m424 < 16; m424 = m424 + 1) 
        begin: inbit424
            assign data_11[m424 + b424*16 + a15*28*16] = data_11_array[a15][b424][m424];
        end
    endgenerate
    generate 
        localparam integer b425 = 5;
        for (m425 = 0; m425 < 16; m425 = m425 + 1) 
        begin: inbit425
            assign data_11[m425 + b425*16 + a15*28*16] = data_11_array[a15][b425][m425];
        end
    endgenerate
    generate 
        localparam integer b426 = 6;
        for (m426 = 0; m426 < 16; m426 = m426 + 1) 
        begin: inbit426
            assign data_11[m426 + b426*16 + a15*28*16] = data_11_array[a15][b426][m426];
        end
    endgenerate
    generate 
        localparam integer b427 = 7;
        for (m427 = 0; m427 < 16; m427 = m427 + 1) 
        begin: inbit427
            assign data_11[m427 + b427*16 + a15*28*16] = data_11_array[a15][b427][m427];
        end
    endgenerate
    generate 
        localparam integer b428 = 8;
        for (m428 = 0; m428 < 16; m428 = m428 + 1) 
        begin: inbit428
            assign data_11[m428 + b428*16 + a15*28*16] = data_11_array[a15][b428][m428];
        end
    endgenerate
    generate 
        localparam integer b429 = 9;
        for (m429 = 0; m429 < 16; m429 = m429 + 1) 
        begin: inbit429
            assign data_11[m429 + b429*16 + a15*28*16] = data_11_array[a15][b429][m429];
        end
    endgenerate
    generate 
        localparam integer b430 = 10;
        for (m430 = 0; m430 < 16; m430 = m430 + 1) 
        begin: inbit430
            assign data_11[m430 + b430*16 + a15*28*16] = data_11_array[a15][b430][m430];
        end
    endgenerate
    generate 
        localparam integer b431 = 11;
        for (m431 = 0; m431 < 16; m431 = m431 + 1) 
        begin: inbit431
            assign data_11[m431 + b431*16 + a15*28*16] = data_11_array[a15][b431][m431];
        end
    endgenerate
    generate 
        localparam integer b432 = 12;
        for (m432 = 0; m432 < 16; m432 = m432 + 1) 
        begin: inbit432
            assign data_11[m432 + b432*16 + a15*28*16] = data_11_array[a15][b432][m432];
        end
    endgenerate
    generate 
        localparam integer b433 = 13;
        for (m433 = 0; m433 < 16; m433 = m433 + 1) 
        begin: inbit433
            assign data_11[m433 + b433*16 + a15*28*16] = data_11_array[a15][b433][m433];
        end
    endgenerate
    generate 
        localparam integer b434 = 14;
        for (m434 = 0; m434 < 16; m434 = m434 + 1) 
        begin: inbit434
            assign data_11[m434 + b434*16 + a15*28*16] = data_11_array[a15][b434][m434];
        end
    endgenerate
    generate 
        localparam integer b435 = 15;
        for (m435 = 0; m435 < 16; m435 = m435 + 1) 
        begin: inbit435
            assign data_11[m435 + b435*16 + a15*28*16] = data_11_array[a15][b435][m435];
        end
    endgenerate
    generate 
        localparam integer b436 = 16;
        for (m436 = 0; m436 < 16; m436 = m436 + 1) 
        begin: inbit436
            assign data_11[m436 + b436*16 + a15*28*16] = data_11_array[a15][b436][m436];
        end
    endgenerate
    generate 
        localparam integer b437 = 17;
        for (m437 = 0; m437 < 16; m437 = m437 + 1) 
        begin: inbit437
            assign data_11[m437 + b437*16 + a15*28*16] = data_11_array[a15][b437][m437];
        end
    endgenerate
    generate 
        localparam integer b438 = 18;
        for (m438 = 0; m438 < 16; m438 = m438 + 1) 
        begin: inbit438
            assign data_11[m438 + b438*16 + a15*28*16] = data_11_array[a15][b438][m438];
        end
    endgenerate
    generate 
        localparam integer b439 = 19;
        for (m439 = 0; m439 < 16; m439 = m439 + 1) 
        begin: inbit439
            assign data_11[m439 + b439*16 + a15*28*16] = data_11_array[a15][b439][m439];
        end
    endgenerate
    generate 
        localparam integer b440 = 20;
        for (m440 = 0; m440 < 16; m440 = m440 + 1) 
        begin: inbit440
            assign data_11[m440 + b440*16 + a15*28*16] = data_11_array[a15][b440][m440];
        end
    endgenerate
    generate 
        localparam integer b441 = 21;
        for (m441 = 0; m441 < 16; m441 = m441 + 1) 
        begin: inbit441
            assign data_11[m441 + b441*16 + a15*28*16] = data_11_array[a15][b441][m441];
        end
    endgenerate
    generate 
        localparam integer b442 = 22;
        for (m442 = 0; m442 < 16; m442 = m442 + 1) 
        begin: inbit442
            assign data_11[m442 + b442*16 + a15*28*16] = data_11_array[a15][b442][m442];
        end
    endgenerate
    generate 
        localparam integer b443 = 23;
        for (m443 = 0; m443 < 16; m443 = m443 + 1) 
        begin: inbit443
            assign data_11[m443 + b443*16 + a15*28*16] = data_11_array[a15][b443][m443];
        end
    endgenerate
    generate 
        localparam integer b444 = 24;
        for (m444 = 0; m444 < 16; m444 = m444 + 1) 
        begin: inbit444
            assign data_11[m444 + b444*16 + a15*28*16] = data_11_array[a15][b444][m444];
        end
    endgenerate
    generate 
        localparam integer b445 = 25;
        for (m445 = 0; m445 < 16; m445 = m445 + 1) 
        begin: inbit445
            assign data_11[m445 + b445*16 + a15*28*16] = data_11_array[a15][b445][m445];
        end
    endgenerate
    generate 
        localparam integer b446 = 26;
        for (m446 = 0; m446 < 16; m446 = m446 + 1) 
        begin: inbit446
            assign data_11[m446 + b446*16 + a15*28*16] = data_11_array[a15][b446][m446];
        end
    endgenerate
    generate 
        localparam integer b447 = 27;
        for (m447 = 0; m447 < 16; m447 = m447 + 1) 
        begin: inbit447
            assign data_11[m447 + b447*16 + a15*28*16] = data_11_array[a15][b447][m447];
        end
    endgenerate
    localparam integer a16 = 16;
    generate 
        localparam integer b448 = 0;
        for (m448 = 0; m448 < 16; m448 = m448 + 1) 
        begin: inbit448
            assign data_11[m448 + b448*16 + a16*28*16] = data_11_array[a16][b448][m448];
        end
    endgenerate
    generate 
        localparam integer b449 = 1;
        for (m449 = 0; m449 < 16; m449 = m449 + 1) 
        begin: inbit449
            assign data_11[m449 + b449*16 + a16*28*16] = data_11_array[a16][b449][m449];
        end
    endgenerate
    generate 
        localparam integer b450 = 2;
        for (m450 = 0; m450 < 16; m450 = m450 + 1) 
        begin: inbit450
            assign data_11[m450 + b450*16 + a16*28*16] = data_11_array[a16][b450][m450];
        end
    endgenerate
    generate 
        localparam integer b451 = 3;
        for (m451 = 0; m451 < 16; m451 = m451 + 1) 
        begin: inbit451
            assign data_11[m451 + b451*16 + a16*28*16] = data_11_array[a16][b451][m451];
        end
    endgenerate
    generate 
        localparam integer b452 = 4;
        for (m452 = 0; m452 < 16; m452 = m452 + 1) 
        begin: inbit452
            assign data_11[m452 + b452*16 + a16*28*16] = data_11_array[a16][b452][m452];
        end
    endgenerate
    generate 
        localparam integer b453 = 5;
        for (m453 = 0; m453 < 16; m453 = m453 + 1) 
        begin: inbit453
            assign data_11[m453 + b453*16 + a16*28*16] = data_11_array[a16][b453][m453];
        end
    endgenerate
    generate 
        localparam integer b454 = 6;
        for (m454 = 0; m454 < 16; m454 = m454 + 1) 
        begin: inbit454
            assign data_11[m454 + b454*16 + a16*28*16] = data_11_array[a16][b454][m454];
        end
    endgenerate
    generate 
        localparam integer b455 = 7;
        for (m455 = 0; m455 < 16; m455 = m455 + 1) 
        begin: inbit455
            assign data_11[m455 + b455*16 + a16*28*16] = data_11_array[a16][b455][m455];
        end
    endgenerate
    generate 
        localparam integer b456 = 8;
        for (m456 = 0; m456 < 16; m456 = m456 + 1) 
        begin: inbit456
            assign data_11[m456 + b456*16 + a16*28*16] = data_11_array[a16][b456][m456];
        end
    endgenerate
    generate 
        localparam integer b457 = 9;
        for (m457 = 0; m457 < 16; m457 = m457 + 1) 
        begin: inbit457
            assign data_11[m457 + b457*16 + a16*28*16] = data_11_array[a16][b457][m457];
        end
    endgenerate
    generate 
        localparam integer b458 = 10;
        for (m458 = 0; m458 < 16; m458 = m458 + 1) 
        begin: inbit458
            assign data_11[m458 + b458*16 + a16*28*16] = data_11_array[a16][b458][m458];
        end
    endgenerate
    generate 
        localparam integer b459 = 11;
        for (m459 = 0; m459 < 16; m459 = m459 + 1) 
        begin: inbit459
            assign data_11[m459 + b459*16 + a16*28*16] = data_11_array[a16][b459][m459];
        end
    endgenerate
    generate 
        localparam integer b460 = 12;
        for (m460 = 0; m460 < 16; m460 = m460 + 1) 
        begin: inbit460
            assign data_11[m460 + b460*16 + a16*28*16] = data_11_array[a16][b460][m460];
        end
    endgenerate
    generate 
        localparam integer b461 = 13;
        for (m461 = 0; m461 < 16; m461 = m461 + 1) 
        begin: inbit461
            assign data_11[m461 + b461*16 + a16*28*16] = data_11_array[a16][b461][m461];
        end
    endgenerate
    generate 
        localparam integer b462 = 14;
        for (m462 = 0; m462 < 16; m462 = m462 + 1) 
        begin: inbit462
            assign data_11[m462 + b462*16 + a16*28*16] = data_11_array[a16][b462][m462];
        end
    endgenerate
    generate 
        localparam integer b463 = 15;
        for (m463 = 0; m463 < 16; m463 = m463 + 1) 
        begin: inbit463
            assign data_11[m463 + b463*16 + a16*28*16] = data_11_array[a16][b463][m463];
        end
    endgenerate
    generate 
        localparam integer b464 = 16;
        for (m464 = 0; m464 < 16; m464 = m464 + 1) 
        begin: inbit464
            assign data_11[m464 + b464*16 + a16*28*16] = data_11_array[a16][b464][m464];
        end
    endgenerate
    generate 
        localparam integer b465 = 17;
        for (m465 = 0; m465 < 16; m465 = m465 + 1) 
        begin: inbit465
            assign data_11[m465 + b465*16 + a16*28*16] = data_11_array[a16][b465][m465];
        end
    endgenerate
    generate 
        localparam integer b466 = 18;
        for (m466 = 0; m466 < 16; m466 = m466 + 1) 
        begin: inbit466
            assign data_11[m466 + b466*16 + a16*28*16] = data_11_array[a16][b466][m466];
        end
    endgenerate
    generate 
        localparam integer b467 = 19;
        for (m467 = 0; m467 < 16; m467 = m467 + 1) 
        begin: inbit467
            assign data_11[m467 + b467*16 + a16*28*16] = data_11_array[a16][b467][m467];
        end
    endgenerate
    generate 
        localparam integer b468 = 20;
        for (m468 = 0; m468 < 16; m468 = m468 + 1) 
        begin: inbit468
            assign data_11[m468 + b468*16 + a16*28*16] = data_11_array[a16][b468][m468];
        end
    endgenerate
    generate 
        localparam integer b469 = 21;
        for (m469 = 0; m469 < 16; m469 = m469 + 1) 
        begin: inbit469
            assign data_11[m469 + b469*16 + a16*28*16] = data_11_array[a16][b469][m469];
        end
    endgenerate
    generate 
        localparam integer b470 = 22;
        for (m470 = 0; m470 < 16; m470 = m470 + 1) 
        begin: inbit470
            assign data_11[m470 + b470*16 + a16*28*16] = data_11_array[a16][b470][m470];
        end
    endgenerate
    generate 
        localparam integer b471 = 23;
        for (m471 = 0; m471 < 16; m471 = m471 + 1) 
        begin: inbit471
            assign data_11[m471 + b471*16 + a16*28*16] = data_11_array[a16][b471][m471];
        end
    endgenerate
    generate 
        localparam integer b472 = 24;
        for (m472 = 0; m472 < 16; m472 = m472 + 1) 
        begin: inbit472
            assign data_11[m472 + b472*16 + a16*28*16] = data_11_array[a16][b472][m472];
        end
    endgenerate
    generate 
        localparam integer b473 = 25;
        for (m473 = 0; m473 < 16; m473 = m473 + 1) 
        begin: inbit473
            assign data_11[m473 + b473*16 + a16*28*16] = data_11_array[a16][b473][m473];
        end
    endgenerate
    generate 
        localparam integer b474 = 26;
        for (m474 = 0; m474 < 16; m474 = m474 + 1) 
        begin: inbit474
            assign data_11[m474 + b474*16 + a16*28*16] = data_11_array[a16][b474][m474];
        end
    endgenerate
    generate 
        localparam integer b475 = 27;
        for (m475 = 0; m475 < 16; m475 = m475 + 1) 
        begin: inbit475
            assign data_11[m475 + b475*16 + a16*28*16] = data_11_array[a16][b475][m475];
        end
    endgenerate
    localparam integer a17 = 17;
    generate 
        localparam integer b476 = 0;
        for (m476 = 0; m476 < 16; m476 = m476 + 1) 
        begin: inbit476
            assign data_11[m476 + b476*16 + a17*28*16] = data_11_array[a17][b476][m476];
        end
    endgenerate
    generate 
        localparam integer b477 = 1;
        for (m477 = 0; m477 < 16; m477 = m477 + 1) 
        begin: inbit477
            assign data_11[m477 + b477*16 + a17*28*16] = data_11_array[a17][b477][m477];
        end
    endgenerate
    generate 
        localparam integer b478 = 2;
        for (m478 = 0; m478 < 16; m478 = m478 + 1) 
        begin: inbit478
            assign data_11[m478 + b478*16 + a17*28*16] = data_11_array[a17][b478][m478];
        end
    endgenerate
    generate 
        localparam integer b479 = 3;
        for (m479 = 0; m479 < 16; m479 = m479 + 1) 
        begin: inbit479
            assign data_11[m479 + b479*16 + a17*28*16] = data_11_array[a17][b479][m479];
        end
    endgenerate
    generate 
        localparam integer b480 = 4;
        for (m480 = 0; m480 < 16; m480 = m480 + 1) 
        begin: inbit480
            assign data_11[m480 + b480*16 + a17*28*16] = data_11_array[a17][b480][m480];
        end
    endgenerate
    generate 
        localparam integer b481 = 5;
        for (m481 = 0; m481 < 16; m481 = m481 + 1) 
        begin: inbit481
            assign data_11[m481 + b481*16 + a17*28*16] = data_11_array[a17][b481][m481];
        end
    endgenerate
    generate 
        localparam integer b482 = 6;
        for (m482 = 0; m482 < 16; m482 = m482 + 1) 
        begin: inbit482
            assign data_11[m482 + b482*16 + a17*28*16] = data_11_array[a17][b482][m482];
        end
    endgenerate
    generate 
        localparam integer b483 = 7;
        for (m483 = 0; m483 < 16; m483 = m483 + 1) 
        begin: inbit483
            assign data_11[m483 + b483*16 + a17*28*16] = data_11_array[a17][b483][m483];
        end
    endgenerate
    generate 
        localparam integer b484 = 8;
        for (m484 = 0; m484 < 16; m484 = m484 + 1) 
        begin: inbit484
            assign data_11[m484 + b484*16 + a17*28*16] = data_11_array[a17][b484][m484];
        end
    endgenerate
    generate 
        localparam integer b485 = 9;
        for (m485 = 0; m485 < 16; m485 = m485 + 1) 
        begin: inbit485
            assign data_11[m485 + b485*16 + a17*28*16] = data_11_array[a17][b485][m485];
        end
    endgenerate
    generate 
        localparam integer b486 = 10;
        for (m486 = 0; m486 < 16; m486 = m486 + 1) 
        begin: inbit486
            assign data_11[m486 + b486*16 + a17*28*16] = data_11_array[a17][b486][m486];
        end
    endgenerate
    generate 
        localparam integer b487 = 11;
        for (m487 = 0; m487 < 16; m487 = m487 + 1) 
        begin: inbit487
            assign data_11[m487 + b487*16 + a17*28*16] = data_11_array[a17][b487][m487];
        end
    endgenerate
    generate 
        localparam integer b488 = 12;
        for (m488 = 0; m488 < 16; m488 = m488 + 1) 
        begin: inbit488
            assign data_11[m488 + b488*16 + a17*28*16] = data_11_array[a17][b488][m488];
        end
    endgenerate
    generate 
        localparam integer b489 = 13;
        for (m489 = 0; m489 < 16; m489 = m489 + 1) 
        begin: inbit489
            assign data_11[m489 + b489*16 + a17*28*16] = data_11_array[a17][b489][m489];
        end
    endgenerate
    generate 
        localparam integer b490 = 14;
        for (m490 = 0; m490 < 16; m490 = m490 + 1) 
        begin: inbit490
            assign data_11[m490 + b490*16 + a17*28*16] = data_11_array[a17][b490][m490];
        end
    endgenerate
    generate 
        localparam integer b491 = 15;
        for (m491 = 0; m491 < 16; m491 = m491 + 1) 
        begin: inbit491
            assign data_11[m491 + b491*16 + a17*28*16] = data_11_array[a17][b491][m491];
        end
    endgenerate
    generate 
        localparam integer b492 = 16;
        for (m492 = 0; m492 < 16; m492 = m492 + 1) 
        begin: inbit492
            assign data_11[m492 + b492*16 + a17*28*16] = data_11_array[a17][b492][m492];
        end
    endgenerate
    generate 
        localparam integer b493 = 17;
        for (m493 = 0; m493 < 16; m493 = m493 + 1) 
        begin: inbit493
            assign data_11[m493 + b493*16 + a17*28*16] = data_11_array[a17][b493][m493];
        end
    endgenerate
    generate 
        localparam integer b494 = 18;
        for (m494 = 0; m494 < 16; m494 = m494 + 1) 
        begin: inbit494
            assign data_11[m494 + b494*16 + a17*28*16] = data_11_array[a17][b494][m494];
        end
    endgenerate
    generate 
        localparam integer b495 = 19;
        for (m495 = 0; m495 < 16; m495 = m495 + 1) 
        begin: inbit495
            assign data_11[m495 + b495*16 + a17*28*16] = data_11_array[a17][b495][m495];
        end
    endgenerate
    generate 
        localparam integer b496 = 20;
        for (m496 = 0; m496 < 16; m496 = m496 + 1) 
        begin: inbit496
            assign data_11[m496 + b496*16 + a17*28*16] = data_11_array[a17][b496][m496];
        end
    endgenerate
    generate 
        localparam integer b497 = 21;
        for (m497 = 0; m497 < 16; m497 = m497 + 1) 
        begin: inbit497
            assign data_11[m497 + b497*16 + a17*28*16] = data_11_array[a17][b497][m497];
        end
    endgenerate
    generate 
        localparam integer b498 = 22;
        for (m498 = 0; m498 < 16; m498 = m498 + 1) 
        begin: inbit498
            assign data_11[m498 + b498*16 + a17*28*16] = data_11_array[a17][b498][m498];
        end
    endgenerate
    generate 
        localparam integer b499 = 23;
        for (m499 = 0; m499 < 16; m499 = m499 + 1) 
        begin: inbit499
            assign data_11[m499 + b499*16 + a17*28*16] = data_11_array[a17][b499][m499];
        end
    endgenerate
    generate 
        localparam integer b500 = 24;
        for (m500 = 0; m500 < 16; m500 = m500 + 1) 
        begin: inbit500
            assign data_11[m500 + b500*16 + a17*28*16] = data_11_array[a17][b500][m500];
        end
    endgenerate
    generate 
        localparam integer b501 = 25;
        for (m501 = 0; m501 < 16; m501 = m501 + 1) 
        begin: inbit501
            assign data_11[m501 + b501*16 + a17*28*16] = data_11_array[a17][b501][m501];
        end
    endgenerate
    generate 
        localparam integer b502 = 26;
        for (m502 = 0; m502 < 16; m502 = m502 + 1) 
        begin: inbit502
            assign data_11[m502 + b502*16 + a17*28*16] = data_11_array[a17][b502][m502];
        end
    endgenerate
    generate 
        localparam integer b503 = 27;
        for (m503 = 0; m503 < 16; m503 = m503 + 1) 
        begin: inbit503
            assign data_11[m503 + b503*16 + a17*28*16] = data_11_array[a17][b503][m503];
        end
    endgenerate
    localparam integer a18 = 18;
    generate 
        localparam integer b504 = 0;
        for (m504 = 0; m504 < 16; m504 = m504 + 1) 
        begin: inbit504
            assign data_11[m504 + b504*16 + a18*28*16] = data_11_array[a18][b504][m504];
        end
    endgenerate
    generate 
        localparam integer b505 = 1;
        for (m505 = 0; m505 < 16; m505 = m505 + 1) 
        begin: inbit505
            assign data_11[m505 + b505*16 + a18*28*16] = data_11_array[a18][b505][m505];
        end
    endgenerate
    generate 
        localparam integer b506 = 2;
        for (m506 = 0; m506 < 16; m506 = m506 + 1) 
        begin: inbit506
            assign data_11[m506 + b506*16 + a18*28*16] = data_11_array[a18][b506][m506];
        end
    endgenerate
    generate 
        localparam integer b507 = 3;
        for (m507 = 0; m507 < 16; m507 = m507 + 1) 
        begin: inbit507
            assign data_11[m507 + b507*16 + a18*28*16] = data_11_array[a18][b507][m507];
        end
    endgenerate
    generate 
        localparam integer b508 = 4;
        for (m508 = 0; m508 < 16; m508 = m508 + 1) 
        begin: inbit508
            assign data_11[m508 + b508*16 + a18*28*16] = data_11_array[a18][b508][m508];
        end
    endgenerate
    generate 
        localparam integer b509 = 5;
        for (m509 = 0; m509 < 16; m509 = m509 + 1) 
        begin: inbit509
            assign data_11[m509 + b509*16 + a18*28*16] = data_11_array[a18][b509][m509];
        end
    endgenerate
    generate 
        localparam integer b510 = 6;
        for (m510 = 0; m510 < 16; m510 = m510 + 1) 
        begin: inbit510
            assign data_11[m510 + b510*16 + a18*28*16] = data_11_array[a18][b510][m510];
        end
    endgenerate
    generate 
        localparam integer b511 = 7;
        for (m511 = 0; m511 < 16; m511 = m511 + 1) 
        begin: inbit511
            assign data_11[m511 + b511*16 + a18*28*16] = data_11_array[a18][b511][m511];
        end
    endgenerate
    generate 
        localparam integer b512 = 8;
        for (m512 = 0; m512 < 16; m512 = m512 + 1) 
        begin: inbit512
            assign data_11[m512 + b512*16 + a18*28*16] = data_11_array[a18][b512][m512];
        end
    endgenerate
    generate 
        localparam integer b513 = 9;
        for (m513 = 0; m513 < 16; m513 = m513 + 1) 
        begin: inbit513
            assign data_11[m513 + b513*16 + a18*28*16] = data_11_array[a18][b513][m513];
        end
    endgenerate
    generate 
        localparam integer b514 = 10;
        for (m514 = 0; m514 < 16; m514 = m514 + 1) 
        begin: inbit514
            assign data_11[m514 + b514*16 + a18*28*16] = data_11_array[a18][b514][m514];
        end
    endgenerate
    generate 
        localparam integer b515 = 11;
        for (m515 = 0; m515 < 16; m515 = m515 + 1) 
        begin: inbit515
            assign data_11[m515 + b515*16 + a18*28*16] = data_11_array[a18][b515][m515];
        end
    endgenerate
    generate 
        localparam integer b516 = 12;
        for (m516 = 0; m516 < 16; m516 = m516 + 1) 
        begin: inbit516
            assign data_11[m516 + b516*16 + a18*28*16] = data_11_array[a18][b516][m516];
        end
    endgenerate
    generate 
        localparam integer b517 = 13;
        for (m517 = 0; m517 < 16; m517 = m517 + 1) 
        begin: inbit517
            assign data_11[m517 + b517*16 + a18*28*16] = data_11_array[a18][b517][m517];
        end
    endgenerate
    generate 
        localparam integer b518 = 14;
        for (m518 = 0; m518 < 16; m518 = m518 + 1) 
        begin: inbit518
            assign data_11[m518 + b518*16 + a18*28*16] = data_11_array[a18][b518][m518];
        end
    endgenerate
    generate 
        localparam integer b519 = 15;
        for (m519 = 0; m519 < 16; m519 = m519 + 1) 
        begin: inbit519
            assign data_11[m519 + b519*16 + a18*28*16] = data_11_array[a18][b519][m519];
        end
    endgenerate
    generate 
        localparam integer b520 = 16;
        for (m520 = 0; m520 < 16; m520 = m520 + 1) 
        begin: inbit520
            assign data_11[m520 + b520*16 + a18*28*16] = data_11_array[a18][b520][m520];
        end
    endgenerate
    generate 
        localparam integer b521 = 17;
        for (m521 = 0; m521 < 16; m521 = m521 + 1) 
        begin: inbit521
            assign data_11[m521 + b521*16 + a18*28*16] = data_11_array[a18][b521][m521];
        end
    endgenerate
    generate 
        localparam integer b522 = 18;
        for (m522 = 0; m522 < 16; m522 = m522 + 1) 
        begin: inbit522
            assign data_11[m522 + b522*16 + a18*28*16] = data_11_array[a18][b522][m522];
        end
    endgenerate
    generate 
        localparam integer b523 = 19;
        for (m523 = 0; m523 < 16; m523 = m523 + 1) 
        begin: inbit523
            assign data_11[m523 + b523*16 + a18*28*16] = data_11_array[a18][b523][m523];
        end
    endgenerate
    generate 
        localparam integer b524 = 20;
        for (m524 = 0; m524 < 16; m524 = m524 + 1) 
        begin: inbit524
            assign data_11[m524 + b524*16 + a18*28*16] = data_11_array[a18][b524][m524];
        end
    endgenerate
    generate 
        localparam integer b525 = 21;
        for (m525 = 0; m525 < 16; m525 = m525 + 1) 
        begin: inbit525
            assign data_11[m525 + b525*16 + a18*28*16] = data_11_array[a18][b525][m525];
        end
    endgenerate
    generate 
        localparam integer b526 = 22;
        for (m526 = 0; m526 < 16; m526 = m526 + 1) 
        begin: inbit526
            assign data_11[m526 + b526*16 + a18*28*16] = data_11_array[a18][b526][m526];
        end
    endgenerate
    generate 
        localparam integer b527 = 23;
        for (m527 = 0; m527 < 16; m527 = m527 + 1) 
        begin: inbit527
            assign data_11[m527 + b527*16 + a18*28*16] = data_11_array[a18][b527][m527];
        end
    endgenerate
    generate 
        localparam integer b528 = 24;
        for (m528 = 0; m528 < 16; m528 = m528 + 1) 
        begin: inbit528
            assign data_11[m528 + b528*16 + a18*28*16] = data_11_array[a18][b528][m528];
        end
    endgenerate
    generate 
        localparam integer b529 = 25;
        for (m529 = 0; m529 < 16; m529 = m529 + 1) 
        begin: inbit529
            assign data_11[m529 + b529*16 + a18*28*16] = data_11_array[a18][b529][m529];
        end
    endgenerate
    generate 
        localparam integer b530 = 26;
        for (m530 = 0; m530 < 16; m530 = m530 + 1) 
        begin: inbit530
            assign data_11[m530 + b530*16 + a18*28*16] = data_11_array[a18][b530][m530];
        end
    endgenerate
    generate 
        localparam integer b531 = 27;
        for (m531 = 0; m531 < 16; m531 = m531 + 1) 
        begin: inbit531
            assign data_11[m531 + b531*16 + a18*28*16] = data_11_array[a18][b531][m531];
        end
    endgenerate
    localparam integer a19 = 19;
    generate 
        localparam integer b532 = 0;
        for (m532 = 0; m532 < 16; m532 = m532 + 1) 
        begin: inbit532
            assign data_11[m532 + b532*16 + a19*28*16] = data_11_array[a19][b532][m532];
        end
    endgenerate
    generate 
        localparam integer b533 = 1;
        for (m533 = 0; m533 < 16; m533 = m533 + 1) 
        begin: inbit533
            assign data_11[m533 + b533*16 + a19*28*16] = data_11_array[a19][b533][m533];
        end
    endgenerate
    generate 
        localparam integer b534 = 2;
        for (m534 = 0; m534 < 16; m534 = m534 + 1) 
        begin: inbit534
            assign data_11[m534 + b534*16 + a19*28*16] = data_11_array[a19][b534][m534];
        end
    endgenerate
    generate 
        localparam integer b535 = 3;
        for (m535 = 0; m535 < 16; m535 = m535 + 1) 
        begin: inbit535
            assign data_11[m535 + b535*16 + a19*28*16] = data_11_array[a19][b535][m535];
        end
    endgenerate
    generate 
        localparam integer b536 = 4;
        for (m536 = 0; m536 < 16; m536 = m536 + 1) 
        begin: inbit536
            assign data_11[m536 + b536*16 + a19*28*16] = data_11_array[a19][b536][m536];
        end
    endgenerate
    generate 
        localparam integer b537 = 5;
        for (m537 = 0; m537 < 16; m537 = m537 + 1) 
        begin: inbit537
            assign data_11[m537 + b537*16 + a19*28*16] = data_11_array[a19][b537][m537];
        end
    endgenerate
    generate 
        localparam integer b538 = 6;
        for (m538 = 0; m538 < 16; m538 = m538 + 1) 
        begin: inbit538
            assign data_11[m538 + b538*16 + a19*28*16] = data_11_array[a19][b538][m538];
        end
    endgenerate
    generate 
        localparam integer b539 = 7;
        for (m539 = 0; m539 < 16; m539 = m539 + 1) 
        begin: inbit539
            assign data_11[m539 + b539*16 + a19*28*16] = data_11_array[a19][b539][m539];
        end
    endgenerate
    generate 
        localparam integer b540 = 8;
        for (m540 = 0; m540 < 16; m540 = m540 + 1) 
        begin: inbit540
            assign data_11[m540 + b540*16 + a19*28*16] = data_11_array[a19][b540][m540];
        end
    endgenerate
    generate 
        localparam integer b541 = 9;
        for (m541 = 0; m541 < 16; m541 = m541 + 1) 
        begin: inbit541
            assign data_11[m541 + b541*16 + a19*28*16] = data_11_array[a19][b541][m541];
        end
    endgenerate
    generate 
        localparam integer b542 = 10;
        for (m542 = 0; m542 < 16; m542 = m542 + 1) 
        begin: inbit542
            assign data_11[m542 + b542*16 + a19*28*16] = data_11_array[a19][b542][m542];
        end
    endgenerate
    generate 
        localparam integer b543 = 11;
        for (m543 = 0; m543 < 16; m543 = m543 + 1) 
        begin: inbit543
            assign data_11[m543 + b543*16 + a19*28*16] = data_11_array[a19][b543][m543];
        end
    endgenerate
    generate 
        localparam integer b544 = 12;
        for (m544 = 0; m544 < 16; m544 = m544 + 1) 
        begin: inbit544
            assign data_11[m544 + b544*16 + a19*28*16] = data_11_array[a19][b544][m544];
        end
    endgenerate
    generate 
        localparam integer b545 = 13;
        for (m545 = 0; m545 < 16; m545 = m545 + 1) 
        begin: inbit545
            assign data_11[m545 + b545*16 + a19*28*16] = data_11_array[a19][b545][m545];
        end
    endgenerate
    generate 
        localparam integer b546 = 14;
        for (m546 = 0; m546 < 16; m546 = m546 + 1) 
        begin: inbit546
            assign data_11[m546 + b546*16 + a19*28*16] = data_11_array[a19][b546][m546];
        end
    endgenerate
    generate 
        localparam integer b547 = 15;
        for (m547 = 0; m547 < 16; m547 = m547 + 1) 
        begin: inbit547
            assign data_11[m547 + b547*16 + a19*28*16] = data_11_array[a19][b547][m547];
        end
    endgenerate
    generate 
        localparam integer b548 = 16;
        for (m548 = 0; m548 < 16; m548 = m548 + 1) 
        begin: inbit548
            assign data_11[m548 + b548*16 + a19*28*16] = data_11_array[a19][b548][m548];
        end
    endgenerate
    generate 
        localparam integer b549 = 17;
        for (m549 = 0; m549 < 16; m549 = m549 + 1) 
        begin: inbit549
            assign data_11[m549 + b549*16 + a19*28*16] = data_11_array[a19][b549][m549];
        end
    endgenerate
    generate 
        localparam integer b550 = 18;
        for (m550 = 0; m550 < 16; m550 = m550 + 1) 
        begin: inbit550
            assign data_11[m550 + b550*16 + a19*28*16] = data_11_array[a19][b550][m550];
        end
    endgenerate
    generate 
        localparam integer b551 = 19;
        for (m551 = 0; m551 < 16; m551 = m551 + 1) 
        begin: inbit551
            assign data_11[m551 + b551*16 + a19*28*16] = data_11_array[a19][b551][m551];
        end
    endgenerate
    generate 
        localparam integer b552 = 20;
        for (m552 = 0; m552 < 16; m552 = m552 + 1) 
        begin: inbit552
            assign data_11[m552 + b552*16 + a19*28*16] = data_11_array[a19][b552][m552];
        end
    endgenerate
    generate 
        localparam integer b553 = 21;
        for (m553 = 0; m553 < 16; m553 = m553 + 1) 
        begin: inbit553
            assign data_11[m553 + b553*16 + a19*28*16] = data_11_array[a19][b553][m553];
        end
    endgenerate
    generate 
        localparam integer b554 = 22;
        for (m554 = 0; m554 < 16; m554 = m554 + 1) 
        begin: inbit554
            assign data_11[m554 + b554*16 + a19*28*16] = data_11_array[a19][b554][m554];
        end
    endgenerate
    generate 
        localparam integer b555 = 23;
        for (m555 = 0; m555 < 16; m555 = m555 + 1) 
        begin: inbit555
            assign data_11[m555 + b555*16 + a19*28*16] = data_11_array[a19][b555][m555];
        end
    endgenerate
    generate 
        localparam integer b556 = 24;
        for (m556 = 0; m556 < 16; m556 = m556 + 1) 
        begin: inbit556
            assign data_11[m556 + b556*16 + a19*28*16] = data_11_array[a19][b556][m556];
        end
    endgenerate
    generate 
        localparam integer b557 = 25;
        for (m557 = 0; m557 < 16; m557 = m557 + 1) 
        begin: inbit557
            assign data_11[m557 + b557*16 + a19*28*16] = data_11_array[a19][b557][m557];
        end
    endgenerate
    generate 
        localparam integer b558 = 26;
        for (m558 = 0; m558 < 16; m558 = m558 + 1) 
        begin: inbit558
            assign data_11[m558 + b558*16 + a19*28*16] = data_11_array[a19][b558][m558];
        end
    endgenerate
    generate 
        localparam integer b559 = 27;
        for (m559 = 0; m559 < 16; m559 = m559 + 1) 
        begin: inbit559
            assign data_11[m559 + b559*16 + a19*28*16] = data_11_array[a19][b559][m559];
        end
    endgenerate
    localparam integer a20 = 20;
    generate 
        localparam integer b560 = 0;
        for (m560 = 0; m560 < 16; m560 = m560 + 1) 
        begin: inbit560
            assign data_11[m560 + b560*16 + a20*28*16] = data_11_array[a20][b560][m560];
        end
    endgenerate
    generate 
        localparam integer b561 = 1;
        for (m561 = 0; m561 < 16; m561 = m561 + 1) 
        begin: inbit561
            assign data_11[m561 + b561*16 + a20*28*16] = data_11_array[a20][b561][m561];
        end
    endgenerate
    generate 
        localparam integer b562 = 2;
        for (m562 = 0; m562 < 16; m562 = m562 + 1) 
        begin: inbit562
            assign data_11[m562 + b562*16 + a20*28*16] = data_11_array[a20][b562][m562];
        end
    endgenerate
    generate 
        localparam integer b563 = 3;
        for (m563 = 0; m563 < 16; m563 = m563 + 1) 
        begin: inbit563
            assign data_11[m563 + b563*16 + a20*28*16] = data_11_array[a20][b563][m563];
        end
    endgenerate
    generate 
        localparam integer b564 = 4;
        for (m564 = 0; m564 < 16; m564 = m564 + 1) 
        begin: inbit564
            assign data_11[m564 + b564*16 + a20*28*16] = data_11_array[a20][b564][m564];
        end
    endgenerate
    generate 
        localparam integer b565 = 5;
        for (m565 = 0; m565 < 16; m565 = m565 + 1) 
        begin: inbit565
            assign data_11[m565 + b565*16 + a20*28*16] = data_11_array[a20][b565][m565];
        end
    endgenerate
    generate 
        localparam integer b566 = 6;
        for (m566 = 0; m566 < 16; m566 = m566 + 1) 
        begin: inbit566
            assign data_11[m566 + b566*16 + a20*28*16] = data_11_array[a20][b566][m566];
        end
    endgenerate
    generate 
        localparam integer b567 = 7;
        for (m567 = 0; m567 < 16; m567 = m567 + 1) 
        begin: inbit567
            assign data_11[m567 + b567*16 + a20*28*16] = data_11_array[a20][b567][m567];
        end
    endgenerate
    generate 
        localparam integer b568 = 8;
        for (m568 = 0; m568 < 16; m568 = m568 + 1) 
        begin: inbit568
            assign data_11[m568 + b568*16 + a20*28*16] = data_11_array[a20][b568][m568];
        end
    endgenerate
    generate 
        localparam integer b569 = 9;
        for (m569 = 0; m569 < 16; m569 = m569 + 1) 
        begin: inbit569
            assign data_11[m569 + b569*16 + a20*28*16] = data_11_array[a20][b569][m569];
        end
    endgenerate
    generate 
        localparam integer b570 = 10;
        for (m570 = 0; m570 < 16; m570 = m570 + 1) 
        begin: inbit570
            assign data_11[m570 + b570*16 + a20*28*16] = data_11_array[a20][b570][m570];
        end
    endgenerate
    generate 
        localparam integer b571 = 11;
        for (m571 = 0; m571 < 16; m571 = m571 + 1) 
        begin: inbit571
            assign data_11[m571 + b571*16 + a20*28*16] = data_11_array[a20][b571][m571];
        end
    endgenerate
    generate 
        localparam integer b572 = 12;
        for (m572 = 0; m572 < 16; m572 = m572 + 1) 
        begin: inbit572
            assign data_11[m572 + b572*16 + a20*28*16] = data_11_array[a20][b572][m572];
        end
    endgenerate
    generate 
        localparam integer b573 = 13;
        for (m573 = 0; m573 < 16; m573 = m573 + 1) 
        begin: inbit573
            assign data_11[m573 + b573*16 + a20*28*16] = data_11_array[a20][b573][m573];
        end
    endgenerate
    generate 
        localparam integer b574 = 14;
        for (m574 = 0; m574 < 16; m574 = m574 + 1) 
        begin: inbit574
            assign data_11[m574 + b574*16 + a20*28*16] = data_11_array[a20][b574][m574];
        end
    endgenerate
    generate 
        localparam integer b575 = 15;
        for (m575 = 0; m575 < 16; m575 = m575 + 1) 
        begin: inbit575
            assign data_11[m575 + b575*16 + a20*28*16] = data_11_array[a20][b575][m575];
        end
    endgenerate
    generate 
        localparam integer b576 = 16;
        for (m576 = 0; m576 < 16; m576 = m576 + 1) 
        begin: inbit576
            assign data_11[m576 + b576*16 + a20*28*16] = data_11_array[a20][b576][m576];
        end
    endgenerate
    generate 
        localparam integer b577 = 17;
        for (m577 = 0; m577 < 16; m577 = m577 + 1) 
        begin: inbit577
            assign data_11[m577 + b577*16 + a20*28*16] = data_11_array[a20][b577][m577];
        end
    endgenerate
    generate 
        localparam integer b578 = 18;
        for (m578 = 0; m578 < 16; m578 = m578 + 1) 
        begin: inbit578
            assign data_11[m578 + b578*16 + a20*28*16] = data_11_array[a20][b578][m578];
        end
    endgenerate
    generate 
        localparam integer b579 = 19;
        for (m579 = 0; m579 < 16; m579 = m579 + 1) 
        begin: inbit579
            assign data_11[m579 + b579*16 + a20*28*16] = data_11_array[a20][b579][m579];
        end
    endgenerate
    generate 
        localparam integer b580 = 20;
        for (m580 = 0; m580 < 16; m580 = m580 + 1) 
        begin: inbit580
            assign data_11[m580 + b580*16 + a20*28*16] = data_11_array[a20][b580][m580];
        end
    endgenerate
    generate 
        localparam integer b581 = 21;
        for (m581 = 0; m581 < 16; m581 = m581 + 1) 
        begin: inbit581
            assign data_11[m581 + b581*16 + a20*28*16] = data_11_array[a20][b581][m581];
        end
    endgenerate
    generate 
        localparam integer b582 = 22;
        for (m582 = 0; m582 < 16; m582 = m582 + 1) 
        begin: inbit582
            assign data_11[m582 + b582*16 + a20*28*16] = data_11_array[a20][b582][m582];
        end
    endgenerate
    generate 
        localparam integer b583 = 23;
        for (m583 = 0; m583 < 16; m583 = m583 + 1) 
        begin: inbit583
            assign data_11[m583 + b583*16 + a20*28*16] = data_11_array[a20][b583][m583];
        end
    endgenerate
    generate 
        localparam integer b584 = 24;
        for (m584 = 0; m584 < 16; m584 = m584 + 1) 
        begin: inbit584
            assign data_11[m584 + b584*16 + a20*28*16] = data_11_array[a20][b584][m584];
        end
    endgenerate
    generate 
        localparam integer b585 = 25;
        for (m585 = 0; m585 < 16; m585 = m585 + 1) 
        begin: inbit585
            assign data_11[m585 + b585*16 + a20*28*16] = data_11_array[a20][b585][m585];
        end
    endgenerate
    generate 
        localparam integer b586 = 26;
        for (m586 = 0; m586 < 16; m586 = m586 + 1) 
        begin: inbit586
            assign data_11[m586 + b586*16 + a20*28*16] = data_11_array[a20][b586][m586];
        end
    endgenerate
    generate 
        localparam integer b587 = 27;
        for (m587 = 0; m587 < 16; m587 = m587 + 1) 
        begin: inbit587
            assign data_11[m587 + b587*16 + a20*28*16] = data_11_array[a20][b587][m587];
        end
    endgenerate
    localparam integer a21 = 21;
    generate 
        localparam integer b588 = 0;
        for (m588 = 0; m588 < 16; m588 = m588 + 1) 
        begin: inbit588
            assign data_11[m588 + b588*16 + a21*28*16] = data_11_array[a21][b588][m588];
        end
    endgenerate
    generate 
        localparam integer b589 = 1;
        for (m589 = 0; m589 < 16; m589 = m589 + 1) 
        begin: inbit589
            assign data_11[m589 + b589*16 + a21*28*16] = data_11_array[a21][b589][m589];
        end
    endgenerate
    generate 
        localparam integer b590 = 2;
        for (m590 = 0; m590 < 16; m590 = m590 + 1) 
        begin: inbit590
            assign data_11[m590 + b590*16 + a21*28*16] = data_11_array[a21][b590][m590];
        end
    endgenerate
    generate 
        localparam integer b591 = 3;
        for (m591 = 0; m591 < 16; m591 = m591 + 1) 
        begin: inbit591
            assign data_11[m591 + b591*16 + a21*28*16] = data_11_array[a21][b591][m591];
        end
    endgenerate
    generate 
        localparam integer b592 = 4;
        for (m592 = 0; m592 < 16; m592 = m592 + 1) 
        begin: inbit592
            assign data_11[m592 + b592*16 + a21*28*16] = data_11_array[a21][b592][m592];
        end
    endgenerate
    generate 
        localparam integer b593 = 5;
        for (m593 = 0; m593 < 16; m593 = m593 + 1) 
        begin: inbit593
            assign data_11[m593 + b593*16 + a21*28*16] = data_11_array[a21][b593][m593];
        end
    endgenerate
    generate 
        localparam integer b594 = 6;
        for (m594 = 0; m594 < 16; m594 = m594 + 1) 
        begin: inbit594
            assign data_11[m594 + b594*16 + a21*28*16] = data_11_array[a21][b594][m594];
        end
    endgenerate
    generate 
        localparam integer b595 = 7;
        for (m595 = 0; m595 < 16; m595 = m595 + 1) 
        begin: inbit595
            assign data_11[m595 + b595*16 + a21*28*16] = data_11_array[a21][b595][m595];
        end
    endgenerate
    generate 
        localparam integer b596 = 8;
        for (m596 = 0; m596 < 16; m596 = m596 + 1) 
        begin: inbit596
            assign data_11[m596 + b596*16 + a21*28*16] = data_11_array[a21][b596][m596];
        end
    endgenerate
    generate 
        localparam integer b597 = 9;
        for (m597 = 0; m597 < 16; m597 = m597 + 1) 
        begin: inbit597
            assign data_11[m597 + b597*16 + a21*28*16] = data_11_array[a21][b597][m597];
        end
    endgenerate
    generate 
        localparam integer b598 = 10;
        for (m598 = 0; m598 < 16; m598 = m598 + 1) 
        begin: inbit598
            assign data_11[m598 + b598*16 + a21*28*16] = data_11_array[a21][b598][m598];
        end
    endgenerate
    generate 
        localparam integer b599 = 11;
        for (m599 = 0; m599 < 16; m599 = m599 + 1) 
        begin: inbit599
            assign data_11[m599 + b599*16 + a21*28*16] = data_11_array[a21][b599][m599];
        end
    endgenerate
    generate 
        localparam integer b600 = 12;
        for (m600 = 0; m600 < 16; m600 = m600 + 1) 
        begin: inbit600
            assign data_11[m600 + b600*16 + a21*28*16] = data_11_array[a21][b600][m600];
        end
    endgenerate
    generate 
        localparam integer b601 = 13;
        for (m601 = 0; m601 < 16; m601 = m601 + 1) 
        begin: inbit601
            assign data_11[m601 + b601*16 + a21*28*16] = data_11_array[a21][b601][m601];
        end
    endgenerate
    generate 
        localparam integer b602 = 14;
        for (m602 = 0; m602 < 16; m602 = m602 + 1) 
        begin: inbit602
            assign data_11[m602 + b602*16 + a21*28*16] = data_11_array[a21][b602][m602];
        end
    endgenerate
    generate 
        localparam integer b603 = 15;
        for (m603 = 0; m603 < 16; m603 = m603 + 1) 
        begin: inbit603
            assign data_11[m603 + b603*16 + a21*28*16] = data_11_array[a21][b603][m603];
        end
    endgenerate
    generate 
        localparam integer b604 = 16;
        for (m604 = 0; m604 < 16; m604 = m604 + 1) 
        begin: inbit604
            assign data_11[m604 + b604*16 + a21*28*16] = data_11_array[a21][b604][m604];
        end
    endgenerate
    generate 
        localparam integer b605 = 17;
        for (m605 = 0; m605 < 16; m605 = m605 + 1) 
        begin: inbit605
            assign data_11[m605 + b605*16 + a21*28*16] = data_11_array[a21][b605][m605];
        end
    endgenerate
    generate 
        localparam integer b606 = 18;
        for (m606 = 0; m606 < 16; m606 = m606 + 1) 
        begin: inbit606
            assign data_11[m606 + b606*16 + a21*28*16] = data_11_array[a21][b606][m606];
        end
    endgenerate
    generate 
        localparam integer b607 = 19;
        for (m607 = 0; m607 < 16; m607 = m607 + 1) 
        begin: inbit607
            assign data_11[m607 + b607*16 + a21*28*16] = data_11_array[a21][b607][m607];
        end
    endgenerate
    generate 
        localparam integer b608 = 20;
        for (m608 = 0; m608 < 16; m608 = m608 + 1) 
        begin: inbit608
            assign data_11[m608 + b608*16 + a21*28*16] = data_11_array[a21][b608][m608];
        end
    endgenerate
    generate 
        localparam integer b609 = 21;
        for (m609 = 0; m609 < 16; m609 = m609 + 1) 
        begin: inbit609
            assign data_11[m609 + b609*16 + a21*28*16] = data_11_array[a21][b609][m609];
        end
    endgenerate
    generate 
        localparam integer b610 = 22;
        for (m610 = 0; m610 < 16; m610 = m610 + 1) 
        begin: inbit610
            assign data_11[m610 + b610*16 + a21*28*16] = data_11_array[a21][b610][m610];
        end
    endgenerate
    generate 
        localparam integer b611 = 23;
        for (m611 = 0; m611 < 16; m611 = m611 + 1) 
        begin: inbit611
            assign data_11[m611 + b611*16 + a21*28*16] = data_11_array[a21][b611][m611];
        end
    endgenerate
    generate 
        localparam integer b612 = 24;
        for (m612 = 0; m612 < 16; m612 = m612 + 1) 
        begin: inbit612
            assign data_11[m612 + b612*16 + a21*28*16] = data_11_array[a21][b612][m612];
        end
    endgenerate
    generate 
        localparam integer b613 = 25;
        for (m613 = 0; m613 < 16; m613 = m613 + 1) 
        begin: inbit613
            assign data_11[m613 + b613*16 + a21*28*16] = data_11_array[a21][b613][m613];
        end
    endgenerate
    generate 
        localparam integer b614 = 26;
        for (m614 = 0; m614 < 16; m614 = m614 + 1) 
        begin: inbit614
            assign data_11[m614 + b614*16 + a21*28*16] = data_11_array[a21][b614][m614];
        end
    endgenerate
    generate 
        localparam integer b615 = 27;
        for (m615 = 0; m615 < 16; m615 = m615 + 1) 
        begin: inbit615
            assign data_11[m615 + b615*16 + a21*28*16] = data_11_array[a21][b615][m615];
        end
    endgenerate
    localparam integer a22 = 22;
    generate 
        localparam integer b616 = 0;
        for (m616 = 0; m616 < 16; m616 = m616 + 1) 
        begin: inbit616
            assign data_11[m616 + b616*16 + a22*28*16] = data_11_array[a22][b616][m616];
        end
    endgenerate
    generate 
        localparam integer b617 = 1;
        for (m617 = 0; m617 < 16; m617 = m617 + 1) 
        begin: inbit617
            assign data_11[m617 + b617*16 + a22*28*16] = data_11_array[a22][b617][m617];
        end
    endgenerate
    generate 
        localparam integer b618 = 2;
        for (m618 = 0; m618 < 16; m618 = m618 + 1) 
        begin: inbit618
            assign data_11[m618 + b618*16 + a22*28*16] = data_11_array[a22][b618][m618];
        end
    endgenerate
    generate 
        localparam integer b619 = 3;
        for (m619 = 0; m619 < 16; m619 = m619 + 1) 
        begin: inbit619
            assign data_11[m619 + b619*16 + a22*28*16] = data_11_array[a22][b619][m619];
        end
    endgenerate
    generate 
        localparam integer b620 = 4;
        for (m620 = 0; m620 < 16; m620 = m620 + 1) 
        begin: inbit620
            assign data_11[m620 + b620*16 + a22*28*16] = data_11_array[a22][b620][m620];
        end
    endgenerate
    generate 
        localparam integer b621 = 5;
        for (m621 = 0; m621 < 16; m621 = m621 + 1) 
        begin: inbit621
            assign data_11[m621 + b621*16 + a22*28*16] = data_11_array[a22][b621][m621];
        end
    endgenerate
    generate 
        localparam integer b622 = 6;
        for (m622 = 0; m622 < 16; m622 = m622 + 1) 
        begin: inbit622
            assign data_11[m622 + b622*16 + a22*28*16] = data_11_array[a22][b622][m622];
        end
    endgenerate
    generate 
        localparam integer b623 = 7;
        for (m623 = 0; m623 < 16; m623 = m623 + 1) 
        begin: inbit623
            assign data_11[m623 + b623*16 + a22*28*16] = data_11_array[a22][b623][m623];
        end
    endgenerate
    generate 
        localparam integer b624 = 8;
        for (m624 = 0; m624 < 16; m624 = m624 + 1) 
        begin: inbit624
            assign data_11[m624 + b624*16 + a22*28*16] = data_11_array[a22][b624][m624];
        end
    endgenerate
    generate 
        localparam integer b625 = 9;
        for (m625 = 0; m625 < 16; m625 = m625 + 1) 
        begin: inbit625
            assign data_11[m625 + b625*16 + a22*28*16] = data_11_array[a22][b625][m625];
        end
    endgenerate
    generate 
        localparam integer b626 = 10;
        for (m626 = 0; m626 < 16; m626 = m626 + 1) 
        begin: inbit626
            assign data_11[m626 + b626*16 + a22*28*16] = data_11_array[a22][b626][m626];
        end
    endgenerate
    generate 
        localparam integer b627 = 11;
        for (m627 = 0; m627 < 16; m627 = m627 + 1) 
        begin: inbit627
            assign data_11[m627 + b627*16 + a22*28*16] = data_11_array[a22][b627][m627];
        end
    endgenerate
    generate 
        localparam integer b628 = 12;
        for (m628 = 0; m628 < 16; m628 = m628 + 1) 
        begin: inbit628
            assign data_11[m628 + b628*16 + a22*28*16] = data_11_array[a22][b628][m628];
        end
    endgenerate
    generate 
        localparam integer b629 = 13;
        for (m629 = 0; m629 < 16; m629 = m629 + 1) 
        begin: inbit629
            assign data_11[m629 + b629*16 + a22*28*16] = data_11_array[a22][b629][m629];
        end
    endgenerate
    generate 
        localparam integer b630 = 14;
        for (m630 = 0; m630 < 16; m630 = m630 + 1) 
        begin: inbit630
            assign data_11[m630 + b630*16 + a22*28*16] = data_11_array[a22][b630][m630];
        end
    endgenerate
    generate 
        localparam integer b631 = 15;
        for (m631 = 0; m631 < 16; m631 = m631 + 1) 
        begin: inbit631
            assign data_11[m631 + b631*16 + a22*28*16] = data_11_array[a22][b631][m631];
        end
    endgenerate
    generate 
        localparam integer b632 = 16;
        for (m632 = 0; m632 < 16; m632 = m632 + 1) 
        begin: inbit632
            assign data_11[m632 + b632*16 + a22*28*16] = data_11_array[a22][b632][m632];
        end
    endgenerate
    generate 
        localparam integer b633 = 17;
        for (m633 = 0; m633 < 16; m633 = m633 + 1) 
        begin: inbit633
            assign data_11[m633 + b633*16 + a22*28*16] = data_11_array[a22][b633][m633];
        end
    endgenerate
    generate 
        localparam integer b634 = 18;
        for (m634 = 0; m634 < 16; m634 = m634 + 1) 
        begin: inbit634
            assign data_11[m634 + b634*16 + a22*28*16] = data_11_array[a22][b634][m634];
        end
    endgenerate
    generate 
        localparam integer b635 = 19;
        for (m635 = 0; m635 < 16; m635 = m635 + 1) 
        begin: inbit635
            assign data_11[m635 + b635*16 + a22*28*16] = data_11_array[a22][b635][m635];
        end
    endgenerate
    generate 
        localparam integer b636 = 20;
        for (m636 = 0; m636 < 16; m636 = m636 + 1) 
        begin: inbit636
            assign data_11[m636 + b636*16 + a22*28*16] = data_11_array[a22][b636][m636];
        end
    endgenerate
    generate 
        localparam integer b637 = 21;
        for (m637 = 0; m637 < 16; m637 = m637 + 1) 
        begin: inbit637
            assign data_11[m637 + b637*16 + a22*28*16] = data_11_array[a22][b637][m637];
        end
    endgenerate
    generate 
        localparam integer b638 = 22;
        for (m638 = 0; m638 < 16; m638 = m638 + 1) 
        begin: inbit638
            assign data_11[m638 + b638*16 + a22*28*16] = data_11_array[a22][b638][m638];
        end
    endgenerate
    generate 
        localparam integer b639 = 23;
        for (m639 = 0; m639 < 16; m639 = m639 + 1) 
        begin: inbit639
            assign data_11[m639 + b639*16 + a22*28*16] = data_11_array[a22][b639][m639];
        end
    endgenerate
    generate 
        localparam integer b640 = 24;
        for (m640 = 0; m640 < 16; m640 = m640 + 1) 
        begin: inbit640
            assign data_11[m640 + b640*16 + a22*28*16] = data_11_array[a22][b640][m640];
        end
    endgenerate
    generate 
        localparam integer b641 = 25;
        for (m641 = 0; m641 < 16; m641 = m641 + 1) 
        begin: inbit641
            assign data_11[m641 + b641*16 + a22*28*16] = data_11_array[a22][b641][m641];
        end
    endgenerate
    generate 
        localparam integer b642 = 26;
        for (m642 = 0; m642 < 16; m642 = m642 + 1) 
        begin: inbit642
            assign data_11[m642 + b642*16 + a22*28*16] = data_11_array[a22][b642][m642];
        end
    endgenerate
    generate 
        localparam integer b643 = 27;
        for (m643 = 0; m643 < 16; m643 = m643 + 1) 
        begin: inbit643
            assign data_11[m643 + b643*16 + a22*28*16] = data_11_array[a22][b643][m643];
        end
    endgenerate
    localparam integer a23 = 23;
    generate 
        localparam integer b644 = 0;
        for (m644 = 0; m644 < 16; m644 = m644 + 1) 
        begin: inbit644
            assign data_11[m644 + b644*16 + a23*28*16] = data_11_array[a23][b644][m644];
        end
    endgenerate
    generate 
        localparam integer b645 = 1;
        for (m645 = 0; m645 < 16; m645 = m645 + 1) 
        begin: inbit645
            assign data_11[m645 + b645*16 + a23*28*16] = data_11_array[a23][b645][m645];
        end
    endgenerate
    generate 
        localparam integer b646 = 2;
        for (m646 = 0; m646 < 16; m646 = m646 + 1) 
        begin: inbit646
            assign data_11[m646 + b646*16 + a23*28*16] = data_11_array[a23][b646][m646];
        end
    endgenerate
    generate 
        localparam integer b647 = 3;
        for (m647 = 0; m647 < 16; m647 = m647 + 1) 
        begin: inbit647
            assign data_11[m647 + b647*16 + a23*28*16] = data_11_array[a23][b647][m647];
        end
    endgenerate
    generate 
        localparam integer b648 = 4;
        for (m648 = 0; m648 < 16; m648 = m648 + 1) 
        begin: inbit648
            assign data_11[m648 + b648*16 + a23*28*16] = data_11_array[a23][b648][m648];
        end
    endgenerate
    generate 
        localparam integer b649 = 5;
        for (m649 = 0; m649 < 16; m649 = m649 + 1) 
        begin: inbit649
            assign data_11[m649 + b649*16 + a23*28*16] = data_11_array[a23][b649][m649];
        end
    endgenerate
    generate 
        localparam integer b650 = 6;
        for (m650 = 0; m650 < 16; m650 = m650 + 1) 
        begin: inbit650
            assign data_11[m650 + b650*16 + a23*28*16] = data_11_array[a23][b650][m650];
        end
    endgenerate
    generate 
        localparam integer b651 = 7;
        for (m651 = 0; m651 < 16; m651 = m651 + 1) 
        begin: inbit651
            assign data_11[m651 + b651*16 + a23*28*16] = data_11_array[a23][b651][m651];
        end
    endgenerate
    generate 
        localparam integer b652 = 8;
        for (m652 = 0; m652 < 16; m652 = m652 + 1) 
        begin: inbit652
            assign data_11[m652 + b652*16 + a23*28*16] = data_11_array[a23][b652][m652];
        end
    endgenerate
    generate 
        localparam integer b653 = 9;
        for (m653 = 0; m653 < 16; m653 = m653 + 1) 
        begin: inbit653
            assign data_11[m653 + b653*16 + a23*28*16] = data_11_array[a23][b653][m653];
        end
    endgenerate
    generate 
        localparam integer b654 = 10;
        for (m654 = 0; m654 < 16; m654 = m654 + 1) 
        begin: inbit654
            assign data_11[m654 + b654*16 + a23*28*16] = data_11_array[a23][b654][m654];
        end
    endgenerate
    generate 
        localparam integer b655 = 11;
        for (m655 = 0; m655 < 16; m655 = m655 + 1) 
        begin: inbit655
            assign data_11[m655 + b655*16 + a23*28*16] = data_11_array[a23][b655][m655];
        end
    endgenerate
    generate 
        localparam integer b656 = 12;
        for (m656 = 0; m656 < 16; m656 = m656 + 1) 
        begin: inbit656
            assign data_11[m656 + b656*16 + a23*28*16] = data_11_array[a23][b656][m656];
        end
    endgenerate
    generate 
        localparam integer b657 = 13;
        for (m657 = 0; m657 < 16; m657 = m657 + 1) 
        begin: inbit657
            assign data_11[m657 + b657*16 + a23*28*16] = data_11_array[a23][b657][m657];
        end
    endgenerate
    generate 
        localparam integer b658 = 14;
        for (m658 = 0; m658 < 16; m658 = m658 + 1) 
        begin: inbit658
            assign data_11[m658 + b658*16 + a23*28*16] = data_11_array[a23][b658][m658];
        end
    endgenerate
    generate 
        localparam integer b659 = 15;
        for (m659 = 0; m659 < 16; m659 = m659 + 1) 
        begin: inbit659
            assign data_11[m659 + b659*16 + a23*28*16] = data_11_array[a23][b659][m659];
        end
    endgenerate
    generate 
        localparam integer b660 = 16;
        for (m660 = 0; m660 < 16; m660 = m660 + 1) 
        begin: inbit660
            assign data_11[m660 + b660*16 + a23*28*16] = data_11_array[a23][b660][m660];
        end
    endgenerate
    generate 
        localparam integer b661 = 17;
        for (m661 = 0; m661 < 16; m661 = m661 + 1) 
        begin: inbit661
            assign data_11[m661 + b661*16 + a23*28*16] = data_11_array[a23][b661][m661];
        end
    endgenerate
    generate 
        localparam integer b662 = 18;
        for (m662 = 0; m662 < 16; m662 = m662 + 1) 
        begin: inbit662
            assign data_11[m662 + b662*16 + a23*28*16] = data_11_array[a23][b662][m662];
        end
    endgenerate
    generate 
        localparam integer b663 = 19;
        for (m663 = 0; m663 < 16; m663 = m663 + 1) 
        begin: inbit663
            assign data_11[m663 + b663*16 + a23*28*16] = data_11_array[a23][b663][m663];
        end
    endgenerate
    generate 
        localparam integer b664 = 20;
        for (m664 = 0; m664 < 16; m664 = m664 + 1) 
        begin: inbit664
            assign data_11[m664 + b664*16 + a23*28*16] = data_11_array[a23][b664][m664];
        end
    endgenerate
    generate 
        localparam integer b665 = 21;
        for (m665 = 0; m665 < 16; m665 = m665 + 1) 
        begin: inbit665
            assign data_11[m665 + b665*16 + a23*28*16] = data_11_array[a23][b665][m665];
        end
    endgenerate
    generate 
        localparam integer b666 = 22;
        for (m666 = 0; m666 < 16; m666 = m666 + 1) 
        begin: inbit666
            assign data_11[m666 + b666*16 + a23*28*16] = data_11_array[a23][b666][m666];
        end
    endgenerate
    generate 
        localparam integer b667 = 23;
        for (m667 = 0; m667 < 16; m667 = m667 + 1) 
        begin: inbit667
            assign data_11[m667 + b667*16 + a23*28*16] = data_11_array[a23][b667][m667];
        end
    endgenerate
    generate 
        localparam integer b668 = 24;
        for (m668 = 0; m668 < 16; m668 = m668 + 1) 
        begin: inbit668
            assign data_11[m668 + b668*16 + a23*28*16] = data_11_array[a23][b668][m668];
        end
    endgenerate
    generate 
        localparam integer b669 = 25;
        for (m669 = 0; m669 < 16; m669 = m669 + 1) 
        begin: inbit669
            assign data_11[m669 + b669*16 + a23*28*16] = data_11_array[a23][b669][m669];
        end
    endgenerate
    generate 
        localparam integer b670 = 26;
        for (m670 = 0; m670 < 16; m670 = m670 + 1) 
        begin: inbit670
            assign data_11[m670 + b670*16 + a23*28*16] = data_11_array[a23][b670][m670];
        end
    endgenerate
    generate 
        localparam integer b671 = 27;
        for (m671 = 0; m671 < 16; m671 = m671 + 1) 
        begin: inbit671
            assign data_11[m671 + b671*16 + a23*28*16] = data_11_array[a23][b671][m671];
        end
    endgenerate
    localparam integer a24 = 24;
    generate 
        localparam integer b672 = 0;
        for (m672 = 0; m672 < 16; m672 = m672 + 1) 
        begin: inbit672
            assign data_11[m672 + b672*16 + a24*28*16] = data_11_array[a24][b672][m672];
        end
    endgenerate
    generate 
        localparam integer b673 = 1;
        for (m673 = 0; m673 < 16; m673 = m673 + 1) 
        begin: inbit673
            assign data_11[m673 + b673*16 + a24*28*16] = data_11_array[a24][b673][m673];
        end
    endgenerate
    generate 
        localparam integer b674 = 2;
        for (m674 = 0; m674 < 16; m674 = m674 + 1) 
        begin: inbit674
            assign data_11[m674 + b674*16 + a24*28*16] = data_11_array[a24][b674][m674];
        end
    endgenerate
    generate 
        localparam integer b675 = 3;
        for (m675 = 0; m675 < 16; m675 = m675 + 1) 
        begin: inbit675
            assign data_11[m675 + b675*16 + a24*28*16] = data_11_array[a24][b675][m675];
        end
    endgenerate
    generate 
        localparam integer b676 = 4;
        for (m676 = 0; m676 < 16; m676 = m676 + 1) 
        begin: inbit676
            assign data_11[m676 + b676*16 + a24*28*16] = data_11_array[a24][b676][m676];
        end
    endgenerate
    generate 
        localparam integer b677 = 5;
        for (m677 = 0; m677 < 16; m677 = m677 + 1) 
        begin: inbit677
            assign data_11[m677 + b677*16 + a24*28*16] = data_11_array[a24][b677][m677];
        end
    endgenerate
    generate 
        localparam integer b678 = 6;
        for (m678 = 0; m678 < 16; m678 = m678 + 1) 
        begin: inbit678
            assign data_11[m678 + b678*16 + a24*28*16] = data_11_array[a24][b678][m678];
        end
    endgenerate
    generate 
        localparam integer b679 = 7;
        for (m679 = 0; m679 < 16; m679 = m679 + 1) 
        begin: inbit679
            assign data_11[m679 + b679*16 + a24*28*16] = data_11_array[a24][b679][m679];
        end
    endgenerate
    generate 
        localparam integer b680 = 8;
        for (m680 = 0; m680 < 16; m680 = m680 + 1) 
        begin: inbit680
            assign data_11[m680 + b680*16 + a24*28*16] = data_11_array[a24][b680][m680];
        end
    endgenerate
    generate 
        localparam integer b681 = 9;
        for (m681 = 0; m681 < 16; m681 = m681 + 1) 
        begin: inbit681
            assign data_11[m681 + b681*16 + a24*28*16] = data_11_array[a24][b681][m681];
        end
    endgenerate
    generate 
        localparam integer b682 = 10;
        for (m682 = 0; m682 < 16; m682 = m682 + 1) 
        begin: inbit682
            assign data_11[m682 + b682*16 + a24*28*16] = data_11_array[a24][b682][m682];
        end
    endgenerate
    generate 
        localparam integer b683 = 11;
        for (m683 = 0; m683 < 16; m683 = m683 + 1) 
        begin: inbit683
            assign data_11[m683 + b683*16 + a24*28*16] = data_11_array[a24][b683][m683];
        end
    endgenerate
    generate 
        localparam integer b684 = 12;
        for (m684 = 0; m684 < 16; m684 = m684 + 1) 
        begin: inbit684
            assign data_11[m684 + b684*16 + a24*28*16] = data_11_array[a24][b684][m684];
        end
    endgenerate
    generate 
        localparam integer b685 = 13;
        for (m685 = 0; m685 < 16; m685 = m685 + 1) 
        begin: inbit685
            assign data_11[m685 + b685*16 + a24*28*16] = data_11_array[a24][b685][m685];
        end
    endgenerate
    generate 
        localparam integer b686 = 14;
        for (m686 = 0; m686 < 16; m686 = m686 + 1) 
        begin: inbit686
            assign data_11[m686 + b686*16 + a24*28*16] = data_11_array[a24][b686][m686];
        end
    endgenerate
    generate 
        localparam integer b687 = 15;
        for (m687 = 0; m687 < 16; m687 = m687 + 1) 
        begin: inbit687
            assign data_11[m687 + b687*16 + a24*28*16] = data_11_array[a24][b687][m687];
        end
    endgenerate
    generate 
        localparam integer b688 = 16;
        for (m688 = 0; m688 < 16; m688 = m688 + 1) 
        begin: inbit688
            assign data_11[m688 + b688*16 + a24*28*16] = data_11_array[a24][b688][m688];
        end
    endgenerate
    generate 
        localparam integer b689 = 17;
        for (m689 = 0; m689 < 16; m689 = m689 + 1) 
        begin: inbit689
            assign data_11[m689 + b689*16 + a24*28*16] = data_11_array[a24][b689][m689];
        end
    endgenerate
    generate 
        localparam integer b690 = 18;
        for (m690 = 0; m690 < 16; m690 = m690 + 1) 
        begin: inbit690
            assign data_11[m690 + b690*16 + a24*28*16] = data_11_array[a24][b690][m690];
        end
    endgenerate
    generate 
        localparam integer b691 = 19;
        for (m691 = 0; m691 < 16; m691 = m691 + 1) 
        begin: inbit691
            assign data_11[m691 + b691*16 + a24*28*16] = data_11_array[a24][b691][m691];
        end
    endgenerate
    generate 
        localparam integer b692 = 20;
        for (m692 = 0; m692 < 16; m692 = m692 + 1) 
        begin: inbit692
            assign data_11[m692 + b692*16 + a24*28*16] = data_11_array[a24][b692][m692];
        end
    endgenerate
    generate 
        localparam integer b693 = 21;
        for (m693 = 0; m693 < 16; m693 = m693 + 1) 
        begin: inbit693
            assign data_11[m693 + b693*16 + a24*28*16] = data_11_array[a24][b693][m693];
        end
    endgenerate
    generate 
        localparam integer b694 = 22;
        for (m694 = 0; m694 < 16; m694 = m694 + 1) 
        begin: inbit694
            assign data_11[m694 + b694*16 + a24*28*16] = data_11_array[a24][b694][m694];
        end
    endgenerate
    generate 
        localparam integer b695 = 23;
        for (m695 = 0; m695 < 16; m695 = m695 + 1) 
        begin: inbit695
            assign data_11[m695 + b695*16 + a24*28*16] = data_11_array[a24][b695][m695];
        end
    endgenerate
    generate 
        localparam integer b696 = 24;
        for (m696 = 0; m696 < 16; m696 = m696 + 1) 
        begin: inbit696
            assign data_11[m696 + b696*16 + a24*28*16] = data_11_array[a24][b696][m696];
        end
    endgenerate
    generate 
        localparam integer b697 = 25;
        for (m697 = 0; m697 < 16; m697 = m697 + 1) 
        begin: inbit697
            assign data_11[m697 + b697*16 + a24*28*16] = data_11_array[a24][b697][m697];
        end
    endgenerate
    generate 
        localparam integer b698 = 26;
        for (m698 = 0; m698 < 16; m698 = m698 + 1) 
        begin: inbit698
            assign data_11[m698 + b698*16 + a24*28*16] = data_11_array[a24][b698][m698];
        end
    endgenerate
    generate 
        localparam integer b699 = 27;
        for (m699 = 0; m699 < 16; m699 = m699 + 1) 
        begin: inbit699
            assign data_11[m699 + b699*16 + a24*28*16] = data_11_array[a24][b699][m699];
        end
    endgenerate
    localparam integer a25 = 25;
    generate 
        localparam integer b700 = 0;
        for (m700 = 0; m700 < 16; m700 = m700 + 1) 
        begin: inbit700
            assign data_11[m700 + b700*16 + a25*28*16] = data_11_array[a25][b700][m700];
        end
    endgenerate
    generate 
        localparam integer b701 = 1;
        for (m701 = 0; m701 < 16; m701 = m701 + 1) 
        begin: inbit701
            assign data_11[m701 + b701*16 + a25*28*16] = data_11_array[a25][b701][m701];
        end
    endgenerate
    generate 
        localparam integer b702 = 2;
        for (m702 = 0; m702 < 16; m702 = m702 + 1) 
        begin: inbit702
            assign data_11[m702 + b702*16 + a25*28*16] = data_11_array[a25][b702][m702];
        end
    endgenerate
    generate 
        localparam integer b703 = 3;
        for (m703 = 0; m703 < 16; m703 = m703 + 1) 
        begin: inbit703
            assign data_11[m703 + b703*16 + a25*28*16] = data_11_array[a25][b703][m703];
        end
    endgenerate
    generate 
        localparam integer b704 = 4;
        for (m704 = 0; m704 < 16; m704 = m704 + 1) 
        begin: inbit704
            assign data_11[m704 + b704*16 + a25*28*16] = data_11_array[a25][b704][m704];
        end
    endgenerate
    generate 
        localparam integer b705 = 5;
        for (m705 = 0; m705 < 16; m705 = m705 + 1) 
        begin: inbit705
            assign data_11[m705 + b705*16 + a25*28*16] = data_11_array[a25][b705][m705];
        end
    endgenerate
    generate 
        localparam integer b706 = 6;
        for (m706 = 0; m706 < 16; m706 = m706 + 1) 
        begin: inbit706
            assign data_11[m706 + b706*16 + a25*28*16] = data_11_array[a25][b706][m706];
        end
    endgenerate
    generate 
        localparam integer b707 = 7;
        for (m707 = 0; m707 < 16; m707 = m707 + 1) 
        begin: inbit707
            assign data_11[m707 + b707*16 + a25*28*16] = data_11_array[a25][b707][m707];
        end
    endgenerate
    generate 
        localparam integer b708 = 8;
        for (m708 = 0; m708 < 16; m708 = m708 + 1) 
        begin: inbit708
            assign data_11[m708 + b708*16 + a25*28*16] = data_11_array[a25][b708][m708];
        end
    endgenerate
    generate 
        localparam integer b709 = 9;
        for (m709 = 0; m709 < 16; m709 = m709 + 1) 
        begin: inbit709
            assign data_11[m709 + b709*16 + a25*28*16] = data_11_array[a25][b709][m709];
        end
    endgenerate
    generate 
        localparam integer b710 = 10;
        for (m710 = 0; m710 < 16; m710 = m710 + 1) 
        begin: inbit710
            assign data_11[m710 + b710*16 + a25*28*16] = data_11_array[a25][b710][m710];
        end
    endgenerate
    generate 
        localparam integer b711 = 11;
        for (m711 = 0; m711 < 16; m711 = m711 + 1) 
        begin: inbit711
            assign data_11[m711 + b711*16 + a25*28*16] = data_11_array[a25][b711][m711];
        end
    endgenerate
    generate 
        localparam integer b712 = 12;
        for (m712 = 0; m712 < 16; m712 = m712 + 1) 
        begin: inbit712
            assign data_11[m712 + b712*16 + a25*28*16] = data_11_array[a25][b712][m712];
        end
    endgenerate
    generate 
        localparam integer b713 = 13;
        for (m713 = 0; m713 < 16; m713 = m713 + 1) 
        begin: inbit713
            assign data_11[m713 + b713*16 + a25*28*16] = data_11_array[a25][b713][m713];
        end
    endgenerate
    generate 
        localparam integer b714 = 14;
        for (m714 = 0; m714 < 16; m714 = m714 + 1) 
        begin: inbit714
            assign data_11[m714 + b714*16 + a25*28*16] = data_11_array[a25][b714][m714];
        end
    endgenerate
    generate 
        localparam integer b715 = 15;
        for (m715 = 0; m715 < 16; m715 = m715 + 1) 
        begin: inbit715
            assign data_11[m715 + b715*16 + a25*28*16] = data_11_array[a25][b715][m715];
        end
    endgenerate
    generate 
        localparam integer b716 = 16;
        for (m716 = 0; m716 < 16; m716 = m716 + 1) 
        begin: inbit716
            assign data_11[m716 + b716*16 + a25*28*16] = data_11_array[a25][b716][m716];
        end
    endgenerate
    generate 
        localparam integer b717 = 17;
        for (m717 = 0; m717 < 16; m717 = m717 + 1) 
        begin: inbit717
            assign data_11[m717 + b717*16 + a25*28*16] = data_11_array[a25][b717][m717];
        end
    endgenerate
    generate 
        localparam integer b718 = 18;
        for (m718 = 0; m718 < 16; m718 = m718 + 1) 
        begin: inbit718
            assign data_11[m718 + b718*16 + a25*28*16] = data_11_array[a25][b718][m718];
        end
    endgenerate
    generate 
        localparam integer b719 = 19;
        for (m719 = 0; m719 < 16; m719 = m719 + 1) 
        begin: inbit719
            assign data_11[m719 + b719*16 + a25*28*16] = data_11_array[a25][b719][m719];
        end
    endgenerate
    generate 
        localparam integer b720 = 20;
        for (m720 = 0; m720 < 16; m720 = m720 + 1) 
        begin: inbit720
            assign data_11[m720 + b720*16 + a25*28*16] = data_11_array[a25][b720][m720];
        end
    endgenerate
    generate 
        localparam integer b721 = 21;
        for (m721 = 0; m721 < 16; m721 = m721 + 1) 
        begin: inbit721
            assign data_11[m721 + b721*16 + a25*28*16] = data_11_array[a25][b721][m721];
        end
    endgenerate
    generate 
        localparam integer b722 = 22;
        for (m722 = 0; m722 < 16; m722 = m722 + 1) 
        begin: inbit722
            assign data_11[m722 + b722*16 + a25*28*16] = data_11_array[a25][b722][m722];
        end
    endgenerate
    generate 
        localparam integer b723 = 23;
        for (m723 = 0; m723 < 16; m723 = m723 + 1) 
        begin: inbit723
            assign data_11[m723 + b723*16 + a25*28*16] = data_11_array[a25][b723][m723];
        end
    endgenerate
    generate 
        localparam integer b724 = 24;
        for (m724 = 0; m724 < 16; m724 = m724 + 1) 
        begin: inbit724
            assign data_11[m724 + b724*16 + a25*28*16] = data_11_array[a25][b724][m724];
        end
    endgenerate
    generate 
        localparam integer b725 = 25;
        for (m725 = 0; m725 < 16; m725 = m725 + 1) 
        begin: inbit725
            assign data_11[m725 + b725*16 + a25*28*16] = data_11_array[a25][b725][m725];
        end
    endgenerate
    generate 
        localparam integer b726 = 26;
        for (m726 = 0; m726 < 16; m726 = m726 + 1) 
        begin: inbit726
            assign data_11[m726 + b726*16 + a25*28*16] = data_11_array[a25][b726][m726];
        end
    endgenerate
    generate 
        localparam integer b727 = 27;
        for (m727 = 0; m727 < 16; m727 = m727 + 1) 
        begin: inbit727
            assign data_11[m727 + b727*16 + a25*28*16] = data_11_array[a25][b727][m727];
        end
    endgenerate
    localparam integer a26 = 26;
    generate 
        localparam integer b728 = 0;
        for (m728 = 0; m728 < 16; m728 = m728 + 1) 
        begin: inbit728
            assign data_11[m728 + b728*16 + a26*28*16] = data_11_array[a26][b728][m728];
        end
    endgenerate
    generate 
        localparam integer b729 = 1;
        for (m729 = 0; m729 < 16; m729 = m729 + 1) 
        begin: inbit729
            assign data_11[m729 + b729*16 + a26*28*16] = data_11_array[a26][b729][m729];
        end
    endgenerate
    generate 
        localparam integer b730 = 2;
        for (m730 = 0; m730 < 16; m730 = m730 + 1) 
        begin: inbit730
            assign data_11[m730 + b730*16 + a26*28*16] = data_11_array[a26][b730][m730];
        end
    endgenerate
    generate 
        localparam integer b731 = 3;
        for (m731 = 0; m731 < 16; m731 = m731 + 1) 
        begin: inbit731
            assign data_11[m731 + b731*16 + a26*28*16] = data_11_array[a26][b731][m731];
        end
    endgenerate
    generate 
        localparam integer b732 = 4;
        for (m732 = 0; m732 < 16; m732 = m732 + 1) 
        begin: inbit732
            assign data_11[m732 + b732*16 + a26*28*16] = data_11_array[a26][b732][m732];
        end
    endgenerate
    generate 
        localparam integer b733 = 5;
        for (m733 = 0; m733 < 16; m733 = m733 + 1) 
        begin: inbit733
            assign data_11[m733 + b733*16 + a26*28*16] = data_11_array[a26][b733][m733];
        end
    endgenerate
    generate 
        localparam integer b734 = 6;
        for (m734 = 0; m734 < 16; m734 = m734 + 1) 
        begin: inbit734
            assign data_11[m734 + b734*16 + a26*28*16] = data_11_array[a26][b734][m734];
        end
    endgenerate
    generate 
        localparam integer b735 = 7;
        for (m735 = 0; m735 < 16; m735 = m735 + 1) 
        begin: inbit735
            assign data_11[m735 + b735*16 + a26*28*16] = data_11_array[a26][b735][m735];
        end
    endgenerate
    generate 
        localparam integer b736 = 8;
        for (m736 = 0; m736 < 16; m736 = m736 + 1) 
        begin: inbit736
            assign data_11[m736 + b736*16 + a26*28*16] = data_11_array[a26][b736][m736];
        end
    endgenerate
    generate 
        localparam integer b737 = 9;
        for (m737 = 0; m737 < 16; m737 = m737 + 1) 
        begin: inbit737
            assign data_11[m737 + b737*16 + a26*28*16] = data_11_array[a26][b737][m737];
        end
    endgenerate
    generate 
        localparam integer b738 = 10;
        for (m738 = 0; m738 < 16; m738 = m738 + 1) 
        begin: inbit738
            assign data_11[m738 + b738*16 + a26*28*16] = data_11_array[a26][b738][m738];
        end
    endgenerate
    generate 
        localparam integer b739 = 11;
        for (m739 = 0; m739 < 16; m739 = m739 + 1) 
        begin: inbit739
            assign data_11[m739 + b739*16 + a26*28*16] = data_11_array[a26][b739][m739];
        end
    endgenerate
    generate 
        localparam integer b740 = 12;
        for (m740 = 0; m740 < 16; m740 = m740 + 1) 
        begin: inbit740
            assign data_11[m740 + b740*16 + a26*28*16] = data_11_array[a26][b740][m740];
        end
    endgenerate
    generate 
        localparam integer b741 = 13;
        for (m741 = 0; m741 < 16; m741 = m741 + 1) 
        begin: inbit741
            assign data_11[m741 + b741*16 + a26*28*16] = data_11_array[a26][b741][m741];
        end
    endgenerate
    generate 
        localparam integer b742 = 14;
        for (m742 = 0; m742 < 16; m742 = m742 + 1) 
        begin: inbit742
            assign data_11[m742 + b742*16 + a26*28*16] = data_11_array[a26][b742][m742];
        end
    endgenerate
    generate 
        localparam integer b743 = 15;
        for (m743 = 0; m743 < 16; m743 = m743 + 1) 
        begin: inbit743
            assign data_11[m743 + b743*16 + a26*28*16] = data_11_array[a26][b743][m743];
        end
    endgenerate
    generate 
        localparam integer b744 = 16;
        for (m744 = 0; m744 < 16; m744 = m744 + 1) 
        begin: inbit744
            assign data_11[m744 + b744*16 + a26*28*16] = data_11_array[a26][b744][m744];
        end
    endgenerate
    generate 
        localparam integer b745 = 17;
        for (m745 = 0; m745 < 16; m745 = m745 + 1) 
        begin: inbit745
            assign data_11[m745 + b745*16 + a26*28*16] = data_11_array[a26][b745][m745];
        end
    endgenerate
    generate 
        localparam integer b746 = 18;
        for (m746 = 0; m746 < 16; m746 = m746 + 1) 
        begin: inbit746
            assign data_11[m746 + b746*16 + a26*28*16] = data_11_array[a26][b746][m746];
        end
    endgenerate
    generate 
        localparam integer b747 = 19;
        for (m747 = 0; m747 < 16; m747 = m747 + 1) 
        begin: inbit747
            assign data_11[m747 + b747*16 + a26*28*16] = data_11_array[a26][b747][m747];
        end
    endgenerate
    generate 
        localparam integer b748 = 20;
        for (m748 = 0; m748 < 16; m748 = m748 + 1) 
        begin: inbit748
            assign data_11[m748 + b748*16 + a26*28*16] = data_11_array[a26][b748][m748];
        end
    endgenerate
    generate 
        localparam integer b749 = 21;
        for (m749 = 0; m749 < 16; m749 = m749 + 1) 
        begin: inbit749
            assign data_11[m749 + b749*16 + a26*28*16] = data_11_array[a26][b749][m749];
        end
    endgenerate
    generate 
        localparam integer b750 = 22;
        for (m750 = 0; m750 < 16; m750 = m750 + 1) 
        begin: inbit750
            assign data_11[m750 + b750*16 + a26*28*16] = data_11_array[a26][b750][m750];
        end
    endgenerate
    generate 
        localparam integer b751 = 23;
        for (m751 = 0; m751 < 16; m751 = m751 + 1) 
        begin: inbit751
            assign data_11[m751 + b751*16 + a26*28*16] = data_11_array[a26][b751][m751];
        end
    endgenerate
    generate 
        localparam integer b752 = 24;
        for (m752 = 0; m752 < 16; m752 = m752 + 1) 
        begin: inbit752
            assign data_11[m752 + b752*16 + a26*28*16] = data_11_array[a26][b752][m752];
        end
    endgenerate
    generate 
        localparam integer b753 = 25;
        for (m753 = 0; m753 < 16; m753 = m753 + 1) 
        begin: inbit753
            assign data_11[m753 + b753*16 + a26*28*16] = data_11_array[a26][b753][m753];
        end
    endgenerate
    generate 
        localparam integer b754 = 26;
        for (m754 = 0; m754 < 16; m754 = m754 + 1) 
        begin: inbit754
            assign data_11[m754 + b754*16 + a26*28*16] = data_11_array[a26][b754][m754];
        end
    endgenerate
    generate 
        localparam integer b755 = 27;
        for (m755 = 0; m755 < 16; m755 = m755 + 1) 
        begin: inbit755
            assign data_11[m755 + b755*16 + a26*28*16] = data_11_array[a26][b755][m755];
        end
    endgenerate
    localparam integer a27 = 27;
    generate 
        localparam integer b756 = 0;
        for (m756 = 0; m756 < 16; m756 = m756 + 1) 
        begin: inbit756
            assign data_11[m756 + b756*16 + a27*28*16] = data_11_array[a27][b756][m756];
        end
    endgenerate
    generate 
        localparam integer b757 = 1;
        for (m757 = 0; m757 < 16; m757 = m757 + 1) 
        begin: inbit757
            assign data_11[m757 + b757*16 + a27*28*16] = data_11_array[a27][b757][m757];
        end
    endgenerate
    generate 
        localparam integer b758 = 2;
        for (m758 = 0; m758 < 16; m758 = m758 + 1) 
        begin: inbit758
            assign data_11[m758 + b758*16 + a27*28*16] = data_11_array[a27][b758][m758];
        end
    endgenerate
    generate 
        localparam integer b759 = 3;
        for (m759 = 0; m759 < 16; m759 = m759 + 1) 
        begin: inbit759
            assign data_11[m759 + b759*16 + a27*28*16] = data_11_array[a27][b759][m759];
        end
    endgenerate
    generate 
        localparam integer b760 = 4;
        for (m760 = 0; m760 < 16; m760 = m760 + 1) 
        begin: inbit760
            assign data_11[m760 + b760*16 + a27*28*16] = data_11_array[a27][b760][m760];
        end
    endgenerate
    generate 
        localparam integer b761 = 5;
        for (m761 = 0; m761 < 16; m761 = m761 + 1) 
        begin: inbit761
            assign data_11[m761 + b761*16 + a27*28*16] = data_11_array[a27][b761][m761];
        end
    endgenerate
    generate 
        localparam integer b762 = 6;
        for (m762 = 0; m762 < 16; m762 = m762 + 1) 
        begin: inbit762
            assign data_11[m762 + b762*16 + a27*28*16] = data_11_array[a27][b762][m762];
        end
    endgenerate
    generate 
        localparam integer b763 = 7;
        for (m763 = 0; m763 < 16; m763 = m763 + 1) 
        begin: inbit763
            assign data_11[m763 + b763*16 + a27*28*16] = data_11_array[a27][b763][m763];
        end
    endgenerate
    generate 
        localparam integer b764 = 8;
        for (m764 = 0; m764 < 16; m764 = m764 + 1) 
        begin: inbit764
            assign data_11[m764 + b764*16 + a27*28*16] = data_11_array[a27][b764][m764];
        end
    endgenerate
    generate 
        localparam integer b765 = 9;
        for (m765 = 0; m765 < 16; m765 = m765 + 1) 
        begin: inbit765
            assign data_11[m765 + b765*16 + a27*28*16] = data_11_array[a27][b765][m765];
        end
    endgenerate
    generate 
        localparam integer b766 = 10;
        for (m766 = 0; m766 < 16; m766 = m766 + 1) 
        begin: inbit766
            assign data_11[m766 + b766*16 + a27*28*16] = data_11_array[a27][b766][m766];
        end
    endgenerate
    generate 
        localparam integer b767 = 11;
        for (m767 = 0; m767 < 16; m767 = m767 + 1) 
        begin: inbit767
            assign data_11[m767 + b767*16 + a27*28*16] = data_11_array[a27][b767][m767];
        end
    endgenerate
    generate 
        localparam integer b768 = 12;
        for (m768 = 0; m768 < 16; m768 = m768 + 1) 
        begin: inbit768
            assign data_11[m768 + b768*16 + a27*28*16] = data_11_array[a27][b768][m768];
        end
    endgenerate
    generate 
        localparam integer b769 = 13;
        for (m769 = 0; m769 < 16; m769 = m769 + 1) 
        begin: inbit769
            assign data_11[m769 + b769*16 + a27*28*16] = data_11_array[a27][b769][m769];
        end
    endgenerate
    generate 
        localparam integer b770 = 14;
        for (m770 = 0; m770 < 16; m770 = m770 + 1) 
        begin: inbit770
            assign data_11[m770 + b770*16 + a27*28*16] = data_11_array[a27][b770][m770];
        end
    endgenerate
    generate 
        localparam integer b771 = 15;
        for (m771 = 0; m771 < 16; m771 = m771 + 1) 
        begin: inbit771
            assign data_11[m771 + b771*16 + a27*28*16] = data_11_array[a27][b771][m771];
        end
    endgenerate
    generate 
        localparam integer b772 = 16;
        for (m772 = 0; m772 < 16; m772 = m772 + 1) 
        begin: inbit772
            assign data_11[m772 + b772*16 + a27*28*16] = data_11_array[a27][b772][m772];
        end
    endgenerate
    generate 
        localparam integer b773 = 17;
        for (m773 = 0; m773 < 16; m773 = m773 + 1) 
        begin: inbit773
            assign data_11[m773 + b773*16 + a27*28*16] = data_11_array[a27][b773][m773];
        end
    endgenerate
    generate 
        localparam integer b774 = 18;
        for (m774 = 0; m774 < 16; m774 = m774 + 1) 
        begin: inbit774
            assign data_11[m774 + b774*16 + a27*28*16] = data_11_array[a27][b774][m774];
        end
    endgenerate
    generate 
        localparam integer b775 = 19;
        for (m775 = 0; m775 < 16; m775 = m775 + 1) 
        begin: inbit775
            assign data_11[m775 + b775*16 + a27*28*16] = data_11_array[a27][b775][m775];
        end
    endgenerate
    generate 
        localparam integer b776 = 20;
        for (m776 = 0; m776 < 16; m776 = m776 + 1) 
        begin: inbit776
            assign data_11[m776 + b776*16 + a27*28*16] = data_11_array[a27][b776][m776];
        end
    endgenerate
    generate 
        localparam integer b777 = 21;
        for (m777 = 0; m777 < 16; m777 = m777 + 1) 
        begin: inbit777
            assign data_11[m777 + b777*16 + a27*28*16] = data_11_array[a27][b777][m777];
        end
    endgenerate
    generate 
        localparam integer b778 = 22;
        for (m778 = 0; m778 < 16; m778 = m778 + 1) 
        begin: inbit778
            assign data_11[m778 + b778*16 + a27*28*16] = data_11_array[a27][b778][m778];
        end
    endgenerate
    generate 
        localparam integer b779 = 23;
        for (m779 = 0; m779 < 16; m779 = m779 + 1) 
        begin: inbit779
            assign data_11[m779 + b779*16 + a27*28*16] = data_11_array[a27][b779][m779];
        end
    endgenerate
    generate 
        localparam integer b780 = 24;
        for (m780 = 0; m780 < 16; m780 = m780 + 1) 
        begin: inbit780
            assign data_11[m780 + b780*16 + a27*28*16] = data_11_array[a27][b780][m780];
        end
    endgenerate
    generate 
        localparam integer b781 = 25;
        for (m781 = 0; m781 < 16; m781 = m781 + 1) 
        begin: inbit781
            assign data_11[m781 + b781*16 + a27*28*16] = data_11_array[a27][b781][m781];
        end
    endgenerate
    generate 
        localparam integer b782 = 26;
        for (m782 = 0; m782 < 16; m782 = m782 + 1) 
        begin: inbit782
            assign data_11[m782 + b782*16 + a27*28*16] = data_11_array[a27][b782][m782];
        end
    endgenerate
    generate 
        localparam integer b783 = 27;
        for (m783 = 0; m783 < 16; m783 = m783 + 1) 
        begin: inbit783
            assign data_11[m783 + b783*16 + a27*28*16] = data_11_array[a27][b783][m783];
        end
    endgenerate
  
  ////ROW 0
  generate
    localparam integer j0 = 0;
    for (i0 = 0; i0 < 24; i0 = i0 + 1)
    begin: addbit0
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j0+0][i0+0]), .Out(multi0[0][i0]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j0+0][i0+1]), .Out(multi0[1][i0]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j0+0][i0+2]), .Out(multi0[2][i0]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j0+0][i0+3]), .Out(multi0[3][i0]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j0+0][i0+4]), .Out(multi0[4][i0]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j0+1][i0+0]), .Out(multi0[5][i0]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j0+1][i0+1]), .Out(multi0[6][i0]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j0+1][i0+2]), .Out(multi0[7][i0]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j0+1][i0+3]), .Out(multi0[8][i0]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j0+1][i0+4]), .Out(multi0[9][i0]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j0+2][i0+0]), .Out(multi0[10][i0]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j0+2][i0+1]), .Out(multi0[11][i0]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j0+2][i0+2]), .Out(multi0[12][i0]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j0+2][i0+3]), .Out(multi0[13][i0]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j0+2][i0+4]), .Out(multi0[14][i0]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j0+3][i0+0]), .Out(multi0[15][i0]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j0+3][i0+1]), .Out(multi0[16][i0]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j0+3][i0+2]), .Out(multi0[17][i0]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j0+3][i0+3]), .Out(multi0[18][i0]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j0+3][i0+4]), .Out(multi0[19][i0]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j0+4][i0+0]), .Out(multi0[20][i0]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j0+4][i0+1]), .Out(multi0[21][i0]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j0+4][i0+2]), .Out(multi0[22][i0]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j0+4][i0+3]), .Out(multi0[23][i0]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j0+4][i0+4]), .Out(multi0[24][i0]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi0[0][i0]), .B(multi0[1][i0]), .Out(sum0[0][i0]));
      FP16_Add stage026(.A(multi0[2][i0]), .B(multi0[3][i0]), .Out(sum0[1][i0]));
      FP16_Add stage027(.A(multi0[4][i0]), .B(multi0[5][i0]), .Out(sum0[2][i0]));
      FP16_Add stage028(.A(multi0[6][i0]), .B(multi0[7][i0]), .Out(sum0[3][i0]));
      FP16_Add stage029(.A(multi0[8][i0]), .B(multi0[9][i0]), .Out(sum0[4][i0]));
      FP16_Add stage030(.A(multi0[10][i0]), .B(multi0[11][i0]), .Out(sum0[5][i0]));
      FP16_Add stage031(.A(multi0[12][i0]), .B(multi0[13][i0]), .Out(sum0[6][i0]));
      FP16_Add stage032(.A(multi0[14][i0]), .B(multi0[15][i0]), .Out(sum0[7][i0]));
      FP16_Add stage033(.A(multi0[16][i0]), .B(multi0[17][i0]), .Out(sum0[8][i0]));
      FP16_Add stage034(.A(multi0[18][i0]), .B(multi0[19][i0]), .Out(sum0[9][i0]));
      FP16_Add stage035(.A(multi0[20][i0]), .B(multi0[21][i0]), .Out(sum0[10][i0]));
      FP16_Add stage036(.A(multi0[22][i0]), .B(multi0[23][i0]), .Out(sum0[11][i0]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum0[0][i0]), .B(sum0[1][i0]), .Out(sum0[12][i0]));
      FP16_Add stage038(.A(sum0[2][i0]), .B(sum0[3][i0]), .Out(sum0[13][i0]));
      FP16_Add stage039(.A(sum0[4][i0]), .B(sum0[5][i0]), .Out(sum0[14][i0]));
      FP16_Add stage040(.A(sum0[6][i0]), .B(sum0[7][i0]), .Out(sum0[15][i0]));
      FP16_Add stage041(.A(sum0[8][i0]), .B(sum0[9][i0]), .Out(sum0[16][i0]));
      FP16_Add stage042(.A(sum0[10][i0]), .B(sum0[11][i0]), .Out(sum0[17][i0]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum0[12][i0]), .B(sum0[13][i0]), .Out(sum0[18][i0]));
      FP16_Add stage044(.A(sum0[14][i0]), .B(sum0[15][i0]), .Out(sum0[19][i0]));
      FP16_Add stage045(.A(sum0[16][i0]), .B(sum0[17][i0]), .Out(sum0[20][i0]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum0[18][i0]), .B(sum0[19][i0]), .Out(sum0[21][i0]));
      FP16_Add stage047(.A(sum0[20][i0]), .B(multi0[24][i0]), .Out(sum0[22][i0]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum0[21][i0]), .B(sum0[22][i0]), .Out(sum0[23][i0]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum0[23][i0]), .B(feature3Bias), .Out(data_11_array[j0][i0]));
    end
  endgenerate
  
  ////ROW 1
  generate
    localparam integer j1 = 1;
    for (i1 = 0; i1 < 24; i1 = i1 + 1)
    begin: addbit1
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j1+0][i1+0]), .Out(multi1[0][i1]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j1+0][i1+1]), .Out(multi1[1][i1]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j1+0][i1+2]), .Out(multi1[2][i1]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j1+0][i1+3]), .Out(multi1[3][i1]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j1+0][i1+4]), .Out(multi1[4][i1]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j1+1][i1+0]), .Out(multi1[5][i1]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j1+1][i1+1]), .Out(multi1[6][i1]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j1+1][i1+2]), .Out(multi1[7][i1]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j1+1][i1+3]), .Out(multi1[8][i1]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j1+1][i1+4]), .Out(multi1[9][i1]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j1+2][i1+0]), .Out(multi1[10][i1]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j1+2][i1+1]), .Out(multi1[11][i1]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j1+2][i1+2]), .Out(multi1[12][i1]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j1+2][i1+3]), .Out(multi1[13][i1]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j1+2][i1+4]), .Out(multi1[14][i1]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j1+3][i1+0]), .Out(multi1[15][i1]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j1+3][i1+1]), .Out(multi1[16][i1]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j1+3][i1+2]), .Out(multi1[17][i1]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j1+3][i1+3]), .Out(multi1[18][i1]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j1+3][i1+4]), .Out(multi1[19][i1]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j1+4][i1+0]), .Out(multi1[20][i1]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j1+4][i1+1]), .Out(multi1[21][i1]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j1+4][i1+2]), .Out(multi1[22][i1]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j1+4][i1+3]), .Out(multi1[23][i1]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j1+4][i1+4]), .Out(multi1[24][i1]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi1[0][i1]), .B(multi1[1][i1]), .Out(sum1[0][i1]));
      FP16_Add stage026(.A(multi1[2][i1]), .B(multi1[3][i1]), .Out(sum1[1][i1]));
      FP16_Add stage027(.A(multi1[4][i1]), .B(multi1[5][i1]), .Out(sum1[2][i1]));
      FP16_Add stage028(.A(multi1[6][i1]), .B(multi1[7][i1]), .Out(sum1[3][i1]));
      FP16_Add stage029(.A(multi1[8][i1]), .B(multi1[9][i1]), .Out(sum1[4][i1]));
      FP16_Add stage030(.A(multi1[10][i1]), .B(multi1[11][i1]), .Out(sum1[5][i1]));
      FP16_Add stage031(.A(multi1[12][i1]), .B(multi1[13][i1]), .Out(sum1[6][i1]));
      FP16_Add stage032(.A(multi1[14][i1]), .B(multi1[15][i1]), .Out(sum1[7][i1]));
      FP16_Add stage033(.A(multi1[16][i1]), .B(multi1[17][i1]), .Out(sum1[8][i1]));
      FP16_Add stage034(.A(multi1[18][i1]), .B(multi1[19][i1]), .Out(sum1[9][i1]));
      FP16_Add stage035(.A(multi1[20][i1]), .B(multi1[21][i1]), .Out(sum1[10][i1]));
      FP16_Add stage036(.A(multi1[22][i1]), .B(multi1[23][i1]), .Out(sum1[11][i1]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum1[0][i1]), .B(sum1[1][i1]), .Out(sum1[12][i1]));
      FP16_Add stage038(.A(sum1[2][i1]), .B(sum1[3][i1]), .Out(sum1[13][i1]));
      FP16_Add stage039(.A(sum1[4][i1]), .B(sum1[5][i1]), .Out(sum1[14][i1]));
      FP16_Add stage040(.A(sum1[6][i1]), .B(sum1[7][i1]), .Out(sum1[15][i1]));
      FP16_Add stage041(.A(sum1[8][i1]), .B(sum1[9][i1]), .Out(sum1[16][i1]));
      FP16_Add stage042(.A(sum1[10][i1]), .B(sum1[11][i1]), .Out(sum1[17][i1]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum1[12][i1]), .B(sum1[13][i1]), .Out(sum1[18][i1]));
      FP16_Add stage044(.A(sum1[14][i1]), .B(sum1[15][i1]), .Out(sum1[19][i1]));
      FP16_Add stage045(.A(sum1[16][i1]), .B(sum1[17][i1]), .Out(sum1[20][i1]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum1[18][i1]), .B(sum1[19][i1]), .Out(sum1[21][i1]));
      FP16_Add stage047(.A(sum1[20][i1]), .B(multi1[24][i1]), .Out(sum1[22][i1]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum1[21][i1]), .B(sum1[22][i1]), .Out(sum1[23][i1]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum1[23][i1]), .B(feature3Bias), .Out(data_11_array[j1][i1]));
    end
  endgenerate
  
  ////ROW 2
  generate
    localparam integer j2 = 2;
    for (i2 = 0; i2 < 24; i2 = i2 + 1)
    begin: addbit2
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j2+0][i2+0]), .Out(multi2[0][i2]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j2+0][i2+1]), .Out(multi2[1][i2]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j2+0][i2+2]), .Out(multi2[2][i2]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j2+0][i2+3]), .Out(multi2[3][i2]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j2+0][i2+4]), .Out(multi2[4][i2]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j2+1][i2+0]), .Out(multi2[5][i2]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j2+1][i2+1]), .Out(multi2[6][i2]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j2+1][i2+2]), .Out(multi2[7][i2]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j2+1][i2+3]), .Out(multi2[8][i2]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j2+1][i2+4]), .Out(multi2[9][i2]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j2+2][i2+0]), .Out(multi2[10][i2]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j2+2][i2+1]), .Out(multi2[11][i2]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j2+2][i2+2]), .Out(multi2[12][i2]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j2+2][i2+3]), .Out(multi2[13][i2]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j2+2][i2+4]), .Out(multi2[14][i2]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j2+3][i2+0]), .Out(multi2[15][i2]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j2+3][i2+1]), .Out(multi2[16][i2]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j2+3][i2+2]), .Out(multi2[17][i2]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j2+3][i2+3]), .Out(multi2[18][i2]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j2+3][i2+4]), .Out(multi2[19][i2]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j2+4][i2+0]), .Out(multi2[20][i2]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j2+4][i2+1]), .Out(multi2[21][i2]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j2+4][i2+2]), .Out(multi2[22][i2]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j2+4][i2+3]), .Out(multi2[23][i2]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j2+4][i2+4]), .Out(multi2[24][i2]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi2[0][i2]), .B(multi2[1][i2]), .Out(sum2[0][i2]));
      FP16_Add stage026(.A(multi2[2][i2]), .B(multi2[3][i2]), .Out(sum2[1][i2]));
      FP16_Add stage027(.A(multi2[4][i2]), .B(multi2[5][i2]), .Out(sum2[2][i2]));
      FP16_Add stage028(.A(multi2[6][i2]), .B(multi2[7][i2]), .Out(sum2[3][i2]));
      FP16_Add stage029(.A(multi2[8][i2]), .B(multi2[9][i2]), .Out(sum2[4][i2]));
      FP16_Add stage030(.A(multi2[10][i2]), .B(multi2[11][i2]), .Out(sum2[5][i2]));
      FP16_Add stage031(.A(multi2[12][i2]), .B(multi2[13][i2]), .Out(sum2[6][i2]));
      FP16_Add stage032(.A(multi2[14][i2]), .B(multi2[15][i2]), .Out(sum2[7][i2]));
      FP16_Add stage033(.A(multi2[16][i2]), .B(multi2[17][i2]), .Out(sum2[8][i2]));
      FP16_Add stage034(.A(multi2[18][i2]), .B(multi2[19][i2]), .Out(sum2[9][i2]));
      FP16_Add stage035(.A(multi2[20][i2]), .B(multi2[21][i2]), .Out(sum2[10][i2]));
      FP16_Add stage036(.A(multi2[22][i2]), .B(multi2[23][i2]), .Out(sum2[11][i2]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum2[0][i2]), .B(sum2[1][i2]), .Out(sum2[12][i2]));
      FP16_Add stage038(.A(sum2[2][i2]), .B(sum2[3][i2]), .Out(sum2[13][i2]));
      FP16_Add stage039(.A(sum2[4][i2]), .B(sum2[5][i2]), .Out(sum2[14][i2]));
      FP16_Add stage040(.A(sum2[6][i2]), .B(sum2[7][i2]), .Out(sum2[15][i2]));
      FP16_Add stage041(.A(sum2[8][i2]), .B(sum2[9][i2]), .Out(sum2[16][i2]));
      FP16_Add stage042(.A(sum2[10][i2]), .B(sum2[11][i2]), .Out(sum2[17][i2]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum2[12][i2]), .B(sum2[13][i2]), .Out(sum2[18][i2]));
      FP16_Add stage044(.A(sum2[14][i2]), .B(sum2[15][i2]), .Out(sum2[19][i2]));
      FP16_Add stage045(.A(sum2[16][i2]), .B(sum2[17][i2]), .Out(sum2[20][i2]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum2[18][i2]), .B(sum2[19][i2]), .Out(sum2[21][i2]));
      FP16_Add stage047(.A(sum2[20][i2]), .B(multi2[24][i2]), .Out(sum2[22][i2]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum2[21][i2]), .B(sum2[22][i2]), .Out(sum2[23][i2]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum2[23][i2]), .B(feature3Bias), .Out(data_11_array[j2][i2]));
    end
  endgenerate
  
  ////ROW 3
  generate
    localparam integer j3 = 3;
    for (i3 = 0; i3 < 24; i3 = i3 + 1)
    begin: addbit3
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j3+0][i3+0]), .Out(multi3[0][i3]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j3+0][i3+1]), .Out(multi3[1][i3]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j3+0][i3+2]), .Out(multi3[2][i3]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j3+0][i3+3]), .Out(multi3[3][i3]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j3+0][i3+4]), .Out(multi3[4][i3]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j3+1][i3+0]), .Out(multi3[5][i3]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j3+1][i3+1]), .Out(multi3[6][i3]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j3+1][i3+2]), .Out(multi3[7][i3]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j3+1][i3+3]), .Out(multi3[8][i3]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j3+1][i3+4]), .Out(multi3[9][i3]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j3+2][i3+0]), .Out(multi3[10][i3]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j3+2][i3+1]), .Out(multi3[11][i3]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j3+2][i3+2]), .Out(multi3[12][i3]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j3+2][i3+3]), .Out(multi3[13][i3]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j3+2][i3+4]), .Out(multi3[14][i3]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j3+3][i3+0]), .Out(multi3[15][i3]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j3+3][i3+1]), .Out(multi3[16][i3]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j3+3][i3+2]), .Out(multi3[17][i3]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j3+3][i3+3]), .Out(multi3[18][i3]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j3+3][i3+4]), .Out(multi3[19][i3]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j3+4][i3+0]), .Out(multi3[20][i3]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j3+4][i3+1]), .Out(multi3[21][i3]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j3+4][i3+2]), .Out(multi3[22][i3]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j3+4][i3+3]), .Out(multi3[23][i3]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j3+4][i3+4]), .Out(multi3[24][i3]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi3[0][i3]), .B(multi3[1][i3]), .Out(sum3[0][i3]));
      FP16_Add stage026(.A(multi3[2][i3]), .B(multi3[3][i3]), .Out(sum3[1][i3]));
      FP16_Add stage027(.A(multi3[4][i3]), .B(multi3[5][i3]), .Out(sum3[2][i3]));
      FP16_Add stage028(.A(multi3[6][i3]), .B(multi3[7][i3]), .Out(sum3[3][i3]));
      FP16_Add stage029(.A(multi3[8][i3]), .B(multi3[9][i3]), .Out(sum3[4][i3]));
      FP16_Add stage030(.A(multi3[10][i3]), .B(multi3[11][i3]), .Out(sum3[5][i3]));
      FP16_Add stage031(.A(multi3[12][i3]), .B(multi3[13][i3]), .Out(sum3[6][i3]));
      FP16_Add stage032(.A(multi3[14][i3]), .B(multi3[15][i3]), .Out(sum3[7][i3]));
      FP16_Add stage033(.A(multi3[16][i3]), .B(multi3[17][i3]), .Out(sum3[8][i3]));
      FP16_Add stage034(.A(multi3[18][i3]), .B(multi3[19][i3]), .Out(sum3[9][i3]));
      FP16_Add stage035(.A(multi3[20][i3]), .B(multi3[21][i3]), .Out(sum3[10][i3]));
      FP16_Add stage036(.A(multi3[22][i3]), .B(multi3[23][i3]), .Out(sum3[11][i3]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum3[0][i3]), .B(sum3[1][i3]), .Out(sum3[12][i3]));
      FP16_Add stage038(.A(sum3[2][i3]), .B(sum3[3][i3]), .Out(sum3[13][i3]));
      FP16_Add stage039(.A(sum3[4][i3]), .B(sum3[5][i3]), .Out(sum3[14][i3]));
      FP16_Add stage040(.A(sum3[6][i3]), .B(sum3[7][i3]), .Out(sum3[15][i3]));
      FP16_Add stage041(.A(sum3[8][i3]), .B(sum3[9][i3]), .Out(sum3[16][i3]));
      FP16_Add stage042(.A(sum3[10][i3]), .B(sum3[11][i3]), .Out(sum3[17][i3]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum3[12][i3]), .B(sum3[13][i3]), .Out(sum3[18][i3]));
      FP16_Add stage044(.A(sum3[14][i3]), .B(sum3[15][i3]), .Out(sum3[19][i3]));
      FP16_Add stage045(.A(sum3[16][i3]), .B(sum3[17][i3]), .Out(sum3[20][i3]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum3[18][i3]), .B(sum3[19][i3]), .Out(sum3[21][i3]));
      FP16_Add stage047(.A(sum3[20][i3]), .B(multi3[24][i3]), .Out(sum3[22][i3]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum3[21][i3]), .B(sum3[22][i3]), .Out(sum3[23][i3]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum3[23][i3]), .B(feature3Bias), .Out(data_11_array[j3][i3]));
    end
  endgenerate
  
  ////ROW 4
  generate
    localparam integer j4 = 4;
    for (i4 = 0; i4 < 24; i4 = i4 + 1)
    begin: addbit4
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j4+0][i4+0]), .Out(multi4[0][i4]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j4+0][i4+1]), .Out(multi4[1][i4]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j4+0][i4+2]), .Out(multi4[2][i4]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j4+0][i4+3]), .Out(multi4[3][i4]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j4+0][i4+4]), .Out(multi4[4][i4]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j4+1][i4+0]), .Out(multi4[5][i4]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j4+1][i4+1]), .Out(multi4[6][i4]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j4+1][i4+2]), .Out(multi4[7][i4]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j4+1][i4+3]), .Out(multi4[8][i4]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j4+1][i4+4]), .Out(multi4[9][i4]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j4+2][i4+0]), .Out(multi4[10][i4]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j4+2][i4+1]), .Out(multi4[11][i4]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j4+2][i4+2]), .Out(multi4[12][i4]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j4+2][i4+3]), .Out(multi4[13][i4]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j4+2][i4+4]), .Out(multi4[14][i4]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j4+3][i4+0]), .Out(multi4[15][i4]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j4+3][i4+1]), .Out(multi4[16][i4]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j4+3][i4+2]), .Out(multi4[17][i4]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j4+3][i4+3]), .Out(multi4[18][i4]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j4+3][i4+4]), .Out(multi4[19][i4]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j4+4][i4+0]), .Out(multi4[20][i4]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j4+4][i4+1]), .Out(multi4[21][i4]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j4+4][i4+2]), .Out(multi4[22][i4]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j4+4][i4+3]), .Out(multi4[23][i4]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j4+4][i4+4]), .Out(multi4[24][i4]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi4[0][i4]), .B(multi4[1][i4]), .Out(sum4[0][i4]));
      FP16_Add stage026(.A(multi4[2][i4]), .B(multi4[3][i4]), .Out(sum4[1][i4]));
      FP16_Add stage027(.A(multi4[4][i4]), .B(multi4[5][i4]), .Out(sum4[2][i4]));
      FP16_Add stage028(.A(multi4[6][i4]), .B(multi4[7][i4]), .Out(sum4[3][i4]));
      FP16_Add stage029(.A(multi4[8][i4]), .B(multi4[9][i4]), .Out(sum4[4][i4]));
      FP16_Add stage030(.A(multi4[10][i4]), .B(multi4[11][i4]), .Out(sum4[5][i4]));
      FP16_Add stage031(.A(multi4[12][i4]), .B(multi4[13][i4]), .Out(sum4[6][i4]));
      FP16_Add stage032(.A(multi4[14][i4]), .B(multi4[15][i4]), .Out(sum4[7][i4]));
      FP16_Add stage033(.A(multi4[16][i4]), .B(multi4[17][i4]), .Out(sum4[8][i4]));
      FP16_Add stage034(.A(multi4[18][i4]), .B(multi4[19][i4]), .Out(sum4[9][i4]));
      FP16_Add stage035(.A(multi4[20][i4]), .B(multi4[21][i4]), .Out(sum4[10][i4]));
      FP16_Add stage036(.A(multi4[22][i4]), .B(multi4[23][i4]), .Out(sum4[11][i4]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum4[0][i4]), .B(sum4[1][i4]), .Out(sum4[12][i4]));
      FP16_Add stage038(.A(sum4[2][i4]), .B(sum4[3][i4]), .Out(sum4[13][i4]));
      FP16_Add stage039(.A(sum4[4][i4]), .B(sum4[5][i4]), .Out(sum4[14][i4]));
      FP16_Add stage040(.A(sum4[6][i4]), .B(sum4[7][i4]), .Out(sum4[15][i4]));
      FP16_Add stage041(.A(sum4[8][i4]), .B(sum4[9][i4]), .Out(sum4[16][i4]));
      FP16_Add stage042(.A(sum4[10][i4]), .B(sum4[11][i4]), .Out(sum4[17][i4]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum4[12][i4]), .B(sum4[13][i4]), .Out(sum4[18][i4]));
      FP16_Add stage044(.A(sum4[14][i4]), .B(sum4[15][i4]), .Out(sum4[19][i4]));
      FP16_Add stage045(.A(sum4[16][i4]), .B(sum4[17][i4]), .Out(sum4[20][i4]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum4[18][i4]), .B(sum4[19][i4]), .Out(sum4[21][i4]));
      FP16_Add stage047(.A(sum4[20][i4]), .B(multi4[24][i4]), .Out(sum4[22][i4]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum4[21][i4]), .B(sum4[22][i4]), .Out(sum4[23][i4]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum4[23][i4]), .B(feature3Bias), .Out(data_11_array[j4][i4]));
    end
  endgenerate
  
  ////ROW 5
  generate
    localparam integer j5 = 5;
    for (i5 = 0; i5 < 24; i5 = i5 + 1)
    begin: addbit5
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j5+0][i5+0]), .Out(multi5[0][i5]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j5+0][i5+1]), .Out(multi5[1][i5]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j5+0][i5+2]), .Out(multi5[2][i5]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j5+0][i5+3]), .Out(multi5[3][i5]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j5+0][i5+4]), .Out(multi5[4][i5]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j5+1][i5+0]), .Out(multi5[5][i5]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j5+1][i5+1]), .Out(multi5[6][i5]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j5+1][i5+2]), .Out(multi5[7][i5]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j5+1][i5+3]), .Out(multi5[8][i5]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j5+1][i5+4]), .Out(multi5[9][i5]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j5+2][i5+0]), .Out(multi5[10][i5]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j5+2][i5+1]), .Out(multi5[11][i5]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j5+2][i5+2]), .Out(multi5[12][i5]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j5+2][i5+3]), .Out(multi5[13][i5]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j5+2][i5+4]), .Out(multi5[14][i5]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j5+3][i5+0]), .Out(multi5[15][i5]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j5+3][i5+1]), .Out(multi5[16][i5]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j5+3][i5+2]), .Out(multi5[17][i5]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j5+3][i5+3]), .Out(multi5[18][i5]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j5+3][i5+4]), .Out(multi5[19][i5]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j5+4][i5+0]), .Out(multi5[20][i5]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j5+4][i5+1]), .Out(multi5[21][i5]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j5+4][i5+2]), .Out(multi5[22][i5]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j5+4][i5+3]), .Out(multi5[23][i5]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j5+4][i5+4]), .Out(multi5[24][i5]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi5[0][i5]), .B(multi5[1][i5]), .Out(sum5[0][i5]));
      FP16_Add stage026(.A(multi5[2][i5]), .B(multi5[3][i5]), .Out(sum5[1][i5]));
      FP16_Add stage027(.A(multi5[4][i5]), .B(multi5[5][i5]), .Out(sum5[2][i5]));
      FP16_Add stage028(.A(multi5[6][i5]), .B(multi5[7][i5]), .Out(sum5[3][i5]));
      FP16_Add stage029(.A(multi5[8][i5]), .B(multi5[9][i5]), .Out(sum5[4][i5]));
      FP16_Add stage030(.A(multi5[10][i5]), .B(multi5[11][i5]), .Out(sum5[5][i5]));
      FP16_Add stage031(.A(multi5[12][i5]), .B(multi5[13][i5]), .Out(sum5[6][i5]));
      FP16_Add stage032(.A(multi5[14][i5]), .B(multi5[15][i5]), .Out(sum5[7][i5]));
      FP16_Add stage033(.A(multi5[16][i5]), .B(multi5[17][i5]), .Out(sum5[8][i5]));
      FP16_Add stage034(.A(multi5[18][i5]), .B(multi5[19][i5]), .Out(sum5[9][i5]));
      FP16_Add stage035(.A(multi5[20][i5]), .B(multi5[21][i5]), .Out(sum5[10][i5]));
      FP16_Add stage036(.A(multi5[22][i5]), .B(multi5[23][i5]), .Out(sum5[11][i5]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum5[0][i5]), .B(sum5[1][i5]), .Out(sum5[12][i5]));
      FP16_Add stage038(.A(sum5[2][i5]), .B(sum5[3][i5]), .Out(sum5[13][i5]));
      FP16_Add stage039(.A(sum5[4][i5]), .B(sum5[5][i5]), .Out(sum5[14][i5]));
      FP16_Add stage040(.A(sum5[6][i5]), .B(sum5[7][i5]), .Out(sum5[15][i5]));
      FP16_Add stage041(.A(sum5[8][i5]), .B(sum5[9][i5]), .Out(sum5[16][i5]));
      FP16_Add stage042(.A(sum5[10][i5]), .B(sum5[11][i5]), .Out(sum5[17][i5]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum5[12][i5]), .B(sum5[13][i5]), .Out(sum5[18][i5]));
      FP16_Add stage044(.A(sum5[14][i5]), .B(sum5[15][i5]), .Out(sum5[19][i5]));
      FP16_Add stage045(.A(sum5[16][i5]), .B(sum5[17][i5]), .Out(sum5[20][i5]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum5[18][i5]), .B(sum5[19][i5]), .Out(sum5[21][i5]));
      FP16_Add stage047(.A(sum5[20][i5]), .B(multi5[24][i5]), .Out(sum5[22][i5]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum5[21][i5]), .B(sum5[22][i5]), .Out(sum5[23][i5]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum5[23][i5]), .B(feature3Bias), .Out(data_11_array[j5][i5]));
    end
  endgenerate
  
  ////ROW 6
  generate
    localparam integer j6 = 6;
    for (i6 = 0; i6 < 24; i6 = i6 + 1)
    begin: addbit6
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j6+0][i6+0]), .Out(multi6[0][i6]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j6+0][i6+1]), .Out(multi6[1][i6]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j6+0][i6+2]), .Out(multi6[2][i6]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j6+0][i6+3]), .Out(multi6[3][i6]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j6+0][i6+4]), .Out(multi6[4][i6]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j6+1][i6+0]), .Out(multi6[5][i6]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j6+1][i6+1]), .Out(multi6[6][i6]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j6+1][i6+2]), .Out(multi6[7][i6]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j6+1][i6+3]), .Out(multi6[8][i6]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j6+1][i6+4]), .Out(multi6[9][i6]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j6+2][i6+0]), .Out(multi6[10][i6]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j6+2][i6+1]), .Out(multi6[11][i6]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j6+2][i6+2]), .Out(multi6[12][i6]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j6+2][i6+3]), .Out(multi6[13][i6]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j6+2][i6+4]), .Out(multi6[14][i6]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j6+3][i6+0]), .Out(multi6[15][i6]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j6+3][i6+1]), .Out(multi6[16][i6]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j6+3][i6+2]), .Out(multi6[17][i6]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j6+3][i6+3]), .Out(multi6[18][i6]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j6+3][i6+4]), .Out(multi6[19][i6]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j6+4][i6+0]), .Out(multi6[20][i6]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j6+4][i6+1]), .Out(multi6[21][i6]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j6+4][i6+2]), .Out(multi6[22][i6]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j6+4][i6+3]), .Out(multi6[23][i6]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j6+4][i6+4]), .Out(multi6[24][i6]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi6[0][i6]), .B(multi6[1][i6]), .Out(sum6[0][i6]));
      FP16_Add stage026(.A(multi6[2][i6]), .B(multi6[3][i6]), .Out(sum6[1][i6]));
      FP16_Add stage027(.A(multi6[4][i6]), .B(multi6[5][i6]), .Out(sum6[2][i6]));
      FP16_Add stage028(.A(multi6[6][i6]), .B(multi6[7][i6]), .Out(sum6[3][i6]));
      FP16_Add stage029(.A(multi6[8][i6]), .B(multi6[9][i6]), .Out(sum6[4][i6]));
      FP16_Add stage030(.A(multi6[10][i6]), .B(multi6[11][i6]), .Out(sum6[5][i6]));
      FP16_Add stage031(.A(multi6[12][i6]), .B(multi6[13][i6]), .Out(sum6[6][i6]));
      FP16_Add stage032(.A(multi6[14][i6]), .B(multi6[15][i6]), .Out(sum6[7][i6]));
      FP16_Add stage033(.A(multi6[16][i6]), .B(multi6[17][i6]), .Out(sum6[8][i6]));
      FP16_Add stage034(.A(multi6[18][i6]), .B(multi6[19][i6]), .Out(sum6[9][i6]));
      FP16_Add stage035(.A(multi6[20][i6]), .B(multi6[21][i6]), .Out(sum6[10][i6]));
      FP16_Add stage036(.A(multi6[22][i6]), .B(multi6[23][i6]), .Out(sum6[11][i6]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum6[0][i6]), .B(sum6[1][i6]), .Out(sum6[12][i6]));
      FP16_Add stage038(.A(sum6[2][i6]), .B(sum6[3][i6]), .Out(sum6[13][i6]));
      FP16_Add stage039(.A(sum6[4][i6]), .B(sum6[5][i6]), .Out(sum6[14][i6]));
      FP16_Add stage040(.A(sum6[6][i6]), .B(sum6[7][i6]), .Out(sum6[15][i6]));
      FP16_Add stage041(.A(sum6[8][i6]), .B(sum6[9][i6]), .Out(sum6[16][i6]));
      FP16_Add stage042(.A(sum6[10][i6]), .B(sum6[11][i6]), .Out(sum6[17][i6]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum6[12][i6]), .B(sum6[13][i6]), .Out(sum6[18][i6]));
      FP16_Add stage044(.A(sum6[14][i6]), .B(sum6[15][i6]), .Out(sum6[19][i6]));
      FP16_Add stage045(.A(sum6[16][i6]), .B(sum6[17][i6]), .Out(sum6[20][i6]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum6[18][i6]), .B(sum6[19][i6]), .Out(sum6[21][i6]));
      FP16_Add stage047(.A(sum6[20][i6]), .B(multi6[24][i6]), .Out(sum6[22][i6]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum6[21][i6]), .B(sum6[22][i6]), .Out(sum6[23][i6]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum6[23][i6]), .B(feature3Bias), .Out(data_11_array[j6][i6]));
    end
  endgenerate
  
  ////ROW 7
  generate
    localparam integer j7 = 7;
    for (i7 = 0; i7 < 24; i7 = i7 + 1)
    begin: addbit7
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j7+0][i7+0]), .Out(multi7[0][i7]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j7+0][i7+1]), .Out(multi7[1][i7]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j7+0][i7+2]), .Out(multi7[2][i7]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j7+0][i7+3]), .Out(multi7[3][i7]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j7+0][i7+4]), .Out(multi7[4][i7]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j7+1][i7+0]), .Out(multi7[5][i7]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j7+1][i7+1]), .Out(multi7[6][i7]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j7+1][i7+2]), .Out(multi7[7][i7]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j7+1][i7+3]), .Out(multi7[8][i7]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j7+1][i7+4]), .Out(multi7[9][i7]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j7+2][i7+0]), .Out(multi7[10][i7]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j7+2][i7+1]), .Out(multi7[11][i7]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j7+2][i7+2]), .Out(multi7[12][i7]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j7+2][i7+3]), .Out(multi7[13][i7]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j7+2][i7+4]), .Out(multi7[14][i7]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j7+3][i7+0]), .Out(multi7[15][i7]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j7+3][i7+1]), .Out(multi7[16][i7]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j7+3][i7+2]), .Out(multi7[17][i7]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j7+3][i7+3]), .Out(multi7[18][i7]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j7+3][i7+4]), .Out(multi7[19][i7]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j7+4][i7+0]), .Out(multi7[20][i7]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j7+4][i7+1]), .Out(multi7[21][i7]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j7+4][i7+2]), .Out(multi7[22][i7]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j7+4][i7+3]), .Out(multi7[23][i7]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j7+4][i7+4]), .Out(multi7[24][i7]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi7[0][i7]), .B(multi7[1][i7]), .Out(sum7[0][i7]));
      FP16_Add stage026(.A(multi7[2][i7]), .B(multi7[3][i7]), .Out(sum7[1][i7]));
      FP16_Add stage027(.A(multi7[4][i7]), .B(multi7[5][i7]), .Out(sum7[2][i7]));
      FP16_Add stage028(.A(multi7[6][i7]), .B(multi7[7][i7]), .Out(sum7[3][i7]));
      FP16_Add stage029(.A(multi7[8][i7]), .B(multi7[9][i7]), .Out(sum7[4][i7]));
      FP16_Add stage030(.A(multi7[10][i7]), .B(multi7[11][i7]), .Out(sum7[5][i7]));
      FP16_Add stage031(.A(multi7[12][i7]), .B(multi7[13][i7]), .Out(sum7[6][i7]));
      FP16_Add stage032(.A(multi7[14][i7]), .B(multi7[15][i7]), .Out(sum7[7][i7]));
      FP16_Add stage033(.A(multi7[16][i7]), .B(multi7[17][i7]), .Out(sum7[8][i7]));
      FP16_Add stage034(.A(multi7[18][i7]), .B(multi7[19][i7]), .Out(sum7[9][i7]));
      FP16_Add stage035(.A(multi7[20][i7]), .B(multi7[21][i7]), .Out(sum7[10][i7]));
      FP16_Add stage036(.A(multi7[22][i7]), .B(multi7[23][i7]), .Out(sum7[11][i7]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum7[0][i7]), .B(sum7[1][i7]), .Out(sum7[12][i7]));
      FP16_Add stage038(.A(sum7[2][i7]), .B(sum7[3][i7]), .Out(sum7[13][i7]));
      FP16_Add stage039(.A(sum7[4][i7]), .B(sum7[5][i7]), .Out(sum7[14][i7]));
      FP16_Add stage040(.A(sum7[6][i7]), .B(sum7[7][i7]), .Out(sum7[15][i7]));
      FP16_Add stage041(.A(sum7[8][i7]), .B(sum7[9][i7]), .Out(sum7[16][i7]));
      FP16_Add stage042(.A(sum7[10][i7]), .B(sum7[11][i7]), .Out(sum7[17][i7]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum7[12][i7]), .B(sum7[13][i7]), .Out(sum7[18][i7]));
      FP16_Add stage044(.A(sum7[14][i7]), .B(sum7[15][i7]), .Out(sum7[19][i7]));
      FP16_Add stage045(.A(sum7[16][i7]), .B(sum7[17][i7]), .Out(sum7[20][i7]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum7[18][i7]), .B(sum7[19][i7]), .Out(sum7[21][i7]));
      FP16_Add stage047(.A(sum7[20][i7]), .B(multi7[24][i7]), .Out(sum7[22][i7]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum7[21][i7]), .B(sum7[22][i7]), .Out(sum7[23][i7]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum7[23][i7]), .B(feature3Bias), .Out(data_11_array[j7][i7]));
    end
  endgenerate
  
  ////ROW 8
  generate
    localparam integer j8 = 8;
    for (i8 = 0; i8 < 24; i8 = i8 + 1)
    begin: addbit8
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j8+0][i8+0]), .Out(multi8[0][i8]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j8+0][i8+1]), .Out(multi8[1][i8]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j8+0][i8+2]), .Out(multi8[2][i8]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j8+0][i8+3]), .Out(multi8[3][i8]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j8+0][i8+4]), .Out(multi8[4][i8]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j8+1][i8+0]), .Out(multi8[5][i8]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j8+1][i8+1]), .Out(multi8[6][i8]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j8+1][i8+2]), .Out(multi8[7][i8]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j8+1][i8+3]), .Out(multi8[8][i8]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j8+1][i8+4]), .Out(multi8[9][i8]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j8+2][i8+0]), .Out(multi8[10][i8]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j8+2][i8+1]), .Out(multi8[11][i8]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j8+2][i8+2]), .Out(multi8[12][i8]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j8+2][i8+3]), .Out(multi8[13][i8]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j8+2][i8+4]), .Out(multi8[14][i8]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j8+3][i8+0]), .Out(multi8[15][i8]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j8+3][i8+1]), .Out(multi8[16][i8]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j8+3][i8+2]), .Out(multi8[17][i8]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j8+3][i8+3]), .Out(multi8[18][i8]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j8+3][i8+4]), .Out(multi8[19][i8]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j8+4][i8+0]), .Out(multi8[20][i8]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j8+4][i8+1]), .Out(multi8[21][i8]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j8+4][i8+2]), .Out(multi8[22][i8]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j8+4][i8+3]), .Out(multi8[23][i8]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j8+4][i8+4]), .Out(multi8[24][i8]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi8[0][i8]), .B(multi8[1][i8]), .Out(sum8[0][i8]));
      FP16_Add stage026(.A(multi8[2][i8]), .B(multi8[3][i8]), .Out(sum8[1][i8]));
      FP16_Add stage027(.A(multi8[4][i8]), .B(multi8[5][i8]), .Out(sum8[2][i8]));
      FP16_Add stage028(.A(multi8[6][i8]), .B(multi8[7][i8]), .Out(sum8[3][i8]));
      FP16_Add stage029(.A(multi8[8][i8]), .B(multi8[9][i8]), .Out(sum8[4][i8]));
      FP16_Add stage030(.A(multi8[10][i8]), .B(multi8[11][i8]), .Out(sum8[5][i8]));
      FP16_Add stage031(.A(multi8[12][i8]), .B(multi8[13][i8]), .Out(sum8[6][i8]));
      FP16_Add stage032(.A(multi8[14][i8]), .B(multi8[15][i8]), .Out(sum8[7][i8]));
      FP16_Add stage033(.A(multi8[16][i8]), .B(multi8[17][i8]), .Out(sum8[8][i8]));
      FP16_Add stage034(.A(multi8[18][i8]), .B(multi8[19][i8]), .Out(sum8[9][i8]));
      FP16_Add stage035(.A(multi8[20][i8]), .B(multi8[21][i8]), .Out(sum8[10][i8]));
      FP16_Add stage036(.A(multi8[22][i8]), .B(multi8[23][i8]), .Out(sum8[11][i8]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum8[0][i8]), .B(sum8[1][i8]), .Out(sum8[12][i8]));
      FP16_Add stage038(.A(sum8[2][i8]), .B(sum8[3][i8]), .Out(sum8[13][i8]));
      FP16_Add stage039(.A(sum8[4][i8]), .B(sum8[5][i8]), .Out(sum8[14][i8]));
      FP16_Add stage040(.A(sum8[6][i8]), .B(sum8[7][i8]), .Out(sum8[15][i8]));
      FP16_Add stage041(.A(sum8[8][i8]), .B(sum8[9][i8]), .Out(sum8[16][i8]));
      FP16_Add stage042(.A(sum8[10][i8]), .B(sum8[11][i8]), .Out(sum8[17][i8]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum8[12][i8]), .B(sum8[13][i8]), .Out(sum8[18][i8]));
      FP16_Add stage044(.A(sum8[14][i8]), .B(sum8[15][i8]), .Out(sum8[19][i8]));
      FP16_Add stage045(.A(sum8[16][i8]), .B(sum8[17][i8]), .Out(sum8[20][i8]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum8[18][i8]), .B(sum8[19][i8]), .Out(sum8[21][i8]));
      FP16_Add stage047(.A(sum8[20][i8]), .B(multi8[24][i8]), .Out(sum8[22][i8]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum8[21][i8]), .B(sum8[22][i8]), .Out(sum8[23][i8]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum8[23][i8]), .B(feature3Bias), .Out(data_11_array[j8][i8]));
    end
  endgenerate
  
  ////ROW 9
  generate
    localparam integer j9 = 9;
    for (i9 = 0; i9 < 24; i9 = i9 + 1)
    begin: addbit9
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j9+0][i9+0]), .Out(multi9[0][i9]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j9+0][i9+1]), .Out(multi9[1][i9]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j9+0][i9+2]), .Out(multi9[2][i9]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j9+0][i9+3]), .Out(multi9[3][i9]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j9+0][i9+4]), .Out(multi9[4][i9]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j9+1][i9+0]), .Out(multi9[5][i9]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j9+1][i9+1]), .Out(multi9[6][i9]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j9+1][i9+2]), .Out(multi9[7][i9]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j9+1][i9+3]), .Out(multi9[8][i9]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j9+1][i9+4]), .Out(multi9[9][i9]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j9+2][i9+0]), .Out(multi9[10][i9]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j9+2][i9+1]), .Out(multi9[11][i9]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j9+2][i9+2]), .Out(multi9[12][i9]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j9+2][i9+3]), .Out(multi9[13][i9]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j9+2][i9+4]), .Out(multi9[14][i9]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j9+3][i9+0]), .Out(multi9[15][i9]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j9+3][i9+1]), .Out(multi9[16][i9]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j9+3][i9+2]), .Out(multi9[17][i9]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j9+3][i9+3]), .Out(multi9[18][i9]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j9+3][i9+4]), .Out(multi9[19][i9]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j9+4][i9+0]), .Out(multi9[20][i9]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j9+4][i9+1]), .Out(multi9[21][i9]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j9+4][i9+2]), .Out(multi9[22][i9]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j9+4][i9+3]), .Out(multi9[23][i9]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j9+4][i9+4]), .Out(multi9[24][i9]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi9[0][i9]), .B(multi9[1][i9]), .Out(sum9[0][i9]));
      FP16_Add stage026(.A(multi9[2][i9]), .B(multi9[3][i9]), .Out(sum9[1][i9]));
      FP16_Add stage027(.A(multi9[4][i9]), .B(multi9[5][i9]), .Out(sum9[2][i9]));
      FP16_Add stage028(.A(multi9[6][i9]), .B(multi9[7][i9]), .Out(sum9[3][i9]));
      FP16_Add stage029(.A(multi9[8][i9]), .B(multi9[9][i9]), .Out(sum9[4][i9]));
      FP16_Add stage030(.A(multi9[10][i9]), .B(multi9[11][i9]), .Out(sum9[5][i9]));
      FP16_Add stage031(.A(multi9[12][i9]), .B(multi9[13][i9]), .Out(sum9[6][i9]));
      FP16_Add stage032(.A(multi9[14][i9]), .B(multi9[15][i9]), .Out(sum9[7][i9]));
      FP16_Add stage033(.A(multi9[16][i9]), .B(multi9[17][i9]), .Out(sum9[8][i9]));
      FP16_Add stage034(.A(multi9[18][i9]), .B(multi9[19][i9]), .Out(sum9[9][i9]));
      FP16_Add stage035(.A(multi9[20][i9]), .B(multi9[21][i9]), .Out(sum9[10][i9]));
      FP16_Add stage036(.A(multi9[22][i9]), .B(multi9[23][i9]), .Out(sum9[11][i9]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum9[0][i9]), .B(sum9[1][i9]), .Out(sum9[12][i9]));
      FP16_Add stage038(.A(sum9[2][i9]), .B(sum9[3][i9]), .Out(sum9[13][i9]));
      FP16_Add stage039(.A(sum9[4][i9]), .B(sum9[5][i9]), .Out(sum9[14][i9]));
      FP16_Add stage040(.A(sum9[6][i9]), .B(sum9[7][i9]), .Out(sum9[15][i9]));
      FP16_Add stage041(.A(sum9[8][i9]), .B(sum9[9][i9]), .Out(sum9[16][i9]));
      FP16_Add stage042(.A(sum9[10][i9]), .B(sum9[11][i9]), .Out(sum9[17][i9]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum9[12][i9]), .B(sum9[13][i9]), .Out(sum9[18][i9]));
      FP16_Add stage044(.A(sum9[14][i9]), .B(sum9[15][i9]), .Out(sum9[19][i9]));
      FP16_Add stage045(.A(sum9[16][i9]), .B(sum9[17][i9]), .Out(sum9[20][i9]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum9[18][i9]), .B(sum9[19][i9]), .Out(sum9[21][i9]));
      FP16_Add stage047(.A(sum9[20][i9]), .B(multi9[24][i9]), .Out(sum9[22][i9]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum9[21][i9]), .B(sum9[22][i9]), .Out(sum9[23][i9]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum9[23][i9]), .B(feature3Bias), .Out(data_11_array[j9][i9]));
    end
  endgenerate
  
  ////ROW 10
  generate
    localparam integer j10 = 10;
    for (i10 = 0; i10 < 24; i10 = i10 + 1)
    begin: addbit10
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j10+0][i10+0]), .Out(multi10[0][i10]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j10+0][i10+1]), .Out(multi10[1][i10]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j10+0][i10+2]), .Out(multi10[2][i10]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j10+0][i10+3]), .Out(multi10[3][i10]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j10+0][i10+4]), .Out(multi10[4][i10]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j10+1][i10+0]), .Out(multi10[5][i10]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j10+1][i10+1]), .Out(multi10[6][i10]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j10+1][i10+2]), .Out(multi10[7][i10]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j10+1][i10+3]), .Out(multi10[8][i10]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j10+1][i10+4]), .Out(multi10[9][i10]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j10+2][i10+0]), .Out(multi10[10][i10]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j10+2][i10+1]), .Out(multi10[11][i10]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j10+2][i10+2]), .Out(multi10[12][i10]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j10+2][i10+3]), .Out(multi10[13][i10]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j10+2][i10+4]), .Out(multi10[14][i10]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j10+3][i10+0]), .Out(multi10[15][i10]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j10+3][i10+1]), .Out(multi10[16][i10]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j10+3][i10+2]), .Out(multi10[17][i10]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j10+3][i10+3]), .Out(multi10[18][i10]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j10+3][i10+4]), .Out(multi10[19][i10]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j10+4][i10+0]), .Out(multi10[20][i10]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j10+4][i10+1]), .Out(multi10[21][i10]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j10+4][i10+2]), .Out(multi10[22][i10]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j10+4][i10+3]), .Out(multi10[23][i10]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j10+4][i10+4]), .Out(multi10[24][i10]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi10[0][i10]), .B(multi10[1][i10]), .Out(sum10[0][i10]));
      FP16_Add stage026(.A(multi10[2][i10]), .B(multi10[3][i10]), .Out(sum10[1][i10]));
      FP16_Add stage027(.A(multi10[4][i10]), .B(multi10[5][i10]), .Out(sum10[2][i10]));
      FP16_Add stage028(.A(multi10[6][i10]), .B(multi10[7][i10]), .Out(sum10[3][i10]));
      FP16_Add stage029(.A(multi10[8][i10]), .B(multi10[9][i10]), .Out(sum10[4][i10]));
      FP16_Add stage030(.A(multi10[10][i10]), .B(multi10[11][i10]), .Out(sum10[5][i10]));
      FP16_Add stage031(.A(multi10[12][i10]), .B(multi10[13][i10]), .Out(sum10[6][i10]));
      FP16_Add stage032(.A(multi10[14][i10]), .B(multi10[15][i10]), .Out(sum10[7][i10]));
      FP16_Add stage033(.A(multi10[16][i10]), .B(multi10[17][i10]), .Out(sum10[8][i10]));
      FP16_Add stage034(.A(multi10[18][i10]), .B(multi10[19][i10]), .Out(sum10[9][i10]));
      FP16_Add stage035(.A(multi10[20][i10]), .B(multi10[21][i10]), .Out(sum10[10][i10]));
      FP16_Add stage036(.A(multi10[22][i10]), .B(multi10[23][i10]), .Out(sum10[11][i10]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum10[0][i10]), .B(sum10[1][i10]), .Out(sum10[12][i10]));
      FP16_Add stage038(.A(sum10[2][i10]), .B(sum10[3][i10]), .Out(sum10[13][i10]));
      FP16_Add stage039(.A(sum10[4][i10]), .B(sum10[5][i10]), .Out(sum10[14][i10]));
      FP16_Add stage040(.A(sum10[6][i10]), .B(sum10[7][i10]), .Out(sum10[15][i10]));
      FP16_Add stage041(.A(sum10[8][i10]), .B(sum10[9][i10]), .Out(sum10[16][i10]));
      FP16_Add stage042(.A(sum10[10][i10]), .B(sum10[11][i10]), .Out(sum10[17][i10]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum10[12][i10]), .B(sum10[13][i10]), .Out(sum10[18][i10]));
      FP16_Add stage044(.A(sum10[14][i10]), .B(sum10[15][i10]), .Out(sum10[19][i10]));
      FP16_Add stage045(.A(sum10[16][i10]), .B(sum10[17][i10]), .Out(sum10[20][i10]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum10[18][i10]), .B(sum10[19][i10]), .Out(sum10[21][i10]));
      FP16_Add stage047(.A(sum10[20][i10]), .B(multi10[24][i10]), .Out(sum10[22][i10]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum10[21][i10]), .B(sum10[22][i10]), .Out(sum10[23][i10]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum10[23][i10]), .B(feature3Bias), .Out(data_11_array[j10][i10]));
    end
  endgenerate
  
    ////ROW 11
  generate
    localparam integer j11 = 11;
    for (i11 = 0; i11 < 24; i11 = i11 + 1)
    begin: addbit11
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j11+0][i11+0]), .Out(multi11[0][i11]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j11+0][i11+1]), .Out(multi11[1][i11]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j11+0][i11+2]), .Out(multi11[2][i11]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j11+0][i11+3]), .Out(multi11[3][i11]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j11+0][i11+4]), .Out(multi11[4][i11]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j11+1][i11+0]), .Out(multi11[5][i11]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j11+1][i11+1]), .Out(multi11[6][i11]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j11+1][i11+2]), .Out(multi11[7][i11]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j11+1][i11+3]), .Out(multi11[8][i11]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j11+1][i11+4]), .Out(multi11[9][i11]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j11+2][i11+0]), .Out(multi11[10][i11]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j11+2][i11+1]), .Out(multi11[11][i11]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j11+2][i11+2]), .Out(multi11[12][i11]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j11+2][i11+3]), .Out(multi11[13][i11]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j11+2][i11+4]), .Out(multi11[14][i11]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j11+3][i11+0]), .Out(multi11[15][i11]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j11+3][i11+1]), .Out(multi11[16][i11]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j11+3][i11+2]), .Out(multi11[17][i11]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j11+3][i11+3]), .Out(multi11[18][i11]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j11+3][i11+4]), .Out(multi11[19][i11]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j11+4][i11+0]), .Out(multi11[20][i11]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j11+4][i11+1]), .Out(multi11[21][i11]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j11+4][i11+2]), .Out(multi11[22][i11]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j11+4][i11+3]), .Out(multi11[23][i11]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j11+4][i11+4]), .Out(multi11[24][i11]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi11[0][i11]), .B(multi11[1][i11]), .Out(sum11[0][i11]));
      FP16_Add stage026(.A(multi11[2][i11]), .B(multi11[3][i11]), .Out(sum11[1][i11]));
      FP16_Add stage027(.A(multi11[4][i11]), .B(multi11[5][i11]), .Out(sum11[2][i11]));
      FP16_Add stage028(.A(multi11[6][i11]), .B(multi11[7][i11]), .Out(sum11[3][i11]));
      FP16_Add stage029(.A(multi11[8][i11]), .B(multi11[9][i11]), .Out(sum11[4][i11]));
      FP16_Add stage030(.A(multi11[10][i11]), .B(multi11[11][i11]), .Out(sum11[5][i11]));
      FP16_Add stage031(.A(multi11[12][i11]), .B(multi11[13][i11]), .Out(sum11[6][i11]));
      FP16_Add stage032(.A(multi11[14][i11]), .B(multi11[15][i11]), .Out(sum11[7][i11]));
      FP16_Add stage033(.A(multi11[16][i11]), .B(multi11[17][i11]), .Out(sum11[8][i11]));
      FP16_Add stage034(.A(multi11[18][i11]), .B(multi11[19][i11]), .Out(sum11[9][i11]));
      FP16_Add stage035(.A(multi11[20][i11]), .B(multi11[21][i11]), .Out(sum11[10][i11]));
      FP16_Add stage036(.A(multi11[22][i11]), .B(multi11[23][i11]), .Out(sum11[11][i11]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum11[0][i11]), .B(sum11[1][i11]), .Out(sum11[12][i11]));
      FP16_Add stage038(.A(sum11[2][i11]), .B(sum11[3][i11]), .Out(sum11[13][i11]));
      FP16_Add stage039(.A(sum11[4][i11]), .B(sum11[5][i11]), .Out(sum11[14][i11]));
      FP16_Add stage040(.A(sum11[6][i11]), .B(sum11[7][i11]), .Out(sum11[15][i11]));
      FP16_Add stage041(.A(sum11[8][i11]), .B(sum11[9][i11]), .Out(sum11[16][i11]));
      FP16_Add stage042(.A(sum11[10][i11]), .B(sum11[11][i11]), .Out(sum11[17][i11]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum11[12][i11]), .B(sum11[13][i11]), .Out(sum11[18][i11]));
      FP16_Add stage044(.A(sum11[14][i11]), .B(sum11[15][i11]), .Out(sum11[19][i11]));
      FP16_Add stage045(.A(sum11[16][i11]), .B(sum11[17][i11]), .Out(sum11[20][i11]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum11[18][i11]), .B(sum11[19][i11]), .Out(sum11[21][i11]));
      FP16_Add stage047(.A(sum11[20][i11]), .B(multi11[24][i11]), .Out(sum11[22][i11]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum11[21][i11]), .B(sum11[22][i11]), .Out(sum11[23][i11]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum11[23][i11]), .B(feature3Bias), .Out(data_11_array[j11][i11]));
    end
  endgenerate

  ////ROW 12
  generate
    localparam integer j12 = 12;
    for (i12 = 0; i12 < 24; i12 = i12 + 1)
    begin: addbit12
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j12+0][i12+0]), .Out(multi12[0][i12]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j12+0][i12+1]), .Out(multi12[1][i12]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j12+0][i12+2]), .Out(multi12[2][i12]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j12+0][i12+3]), .Out(multi12[3][i12]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j12+0][i12+4]), .Out(multi12[4][i12]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j12+1][i12+0]), .Out(multi12[5][i12]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j12+1][i12+1]), .Out(multi12[6][i12]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j12+1][i12+2]), .Out(multi12[7][i12]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j12+1][i12+3]), .Out(multi12[8][i12]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j12+1][i12+4]), .Out(multi12[9][i12]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j12+2][i12+0]), .Out(multi12[10][i12]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j12+2][i12+1]), .Out(multi12[11][i12]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j12+2][i12+2]), .Out(multi12[12][i12]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j12+2][i12+3]), .Out(multi12[13][i12]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j12+2][i12+4]), .Out(multi12[14][i12]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j12+3][i12+0]), .Out(multi12[15][i12]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j12+3][i12+1]), .Out(multi12[16][i12]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j12+3][i12+2]), .Out(multi12[17][i12]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j12+3][i12+3]), .Out(multi12[18][i12]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j12+3][i12+4]), .Out(multi12[19][i12]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j12+4][i12+0]), .Out(multi12[20][i12]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j12+4][i12+1]), .Out(multi12[21][i12]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j12+4][i12+2]), .Out(multi12[22][i12]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j12+4][i12+3]), .Out(multi12[23][i12]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j12+4][i12+4]), .Out(multi12[24][i12]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi12[0][i12]), .B(multi12[1][i12]), .Out(sum12[0][i12]));
      FP16_Add stage026(.A(multi12[2][i12]), .B(multi12[3][i12]), .Out(sum12[1][i12]));
      FP16_Add stage027(.A(multi12[4][i12]), .B(multi12[5][i12]), .Out(sum12[2][i12]));
      FP16_Add stage028(.A(multi12[6][i12]), .B(multi12[7][i12]), .Out(sum12[3][i12]));
      FP16_Add stage029(.A(multi12[8][i12]), .B(multi12[9][i12]), .Out(sum12[4][i12]));
      FP16_Add stage030(.A(multi12[10][i12]), .B(multi12[11][i12]), .Out(sum12[5][i12]));
      FP16_Add stage031(.A(multi12[12][i12]), .B(multi12[13][i12]), .Out(sum12[6][i12]));
      FP16_Add stage032(.A(multi12[14][i12]), .B(multi12[15][i12]), .Out(sum12[7][i12]));
      FP16_Add stage033(.A(multi12[16][i12]), .B(multi12[17][i12]), .Out(sum12[8][i12]));
      FP16_Add stage034(.A(multi12[18][i12]), .B(multi12[19][i12]), .Out(sum12[9][i12]));
      FP16_Add stage035(.A(multi12[20][i12]), .B(multi12[21][i12]), .Out(sum12[10][i12]));
      FP16_Add stage036(.A(multi12[22][i12]), .B(multi12[23][i12]), .Out(sum12[11][i12]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum12[0][i12]), .B(sum12[1][i12]), .Out(sum12[12][i12]));
      FP16_Add stage038(.A(sum12[2][i12]), .B(sum12[3][i12]), .Out(sum12[13][i12]));
      FP16_Add stage039(.A(sum12[4][i12]), .B(sum12[5][i12]), .Out(sum12[14][i12]));
      FP16_Add stage040(.A(sum12[6][i12]), .B(sum12[7][i12]), .Out(sum12[15][i12]));
      FP16_Add stage041(.A(sum12[8][i12]), .B(sum12[9][i12]), .Out(sum12[16][i12]));
      FP16_Add stage042(.A(sum12[10][i12]), .B(sum12[11][i12]), .Out(sum12[17][i12]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum12[12][i12]), .B(sum12[13][i12]), .Out(sum12[18][i12]));
      FP16_Add stage044(.A(sum12[14][i12]), .B(sum12[15][i12]), .Out(sum12[19][i12]));
      FP16_Add stage045(.A(sum12[16][i12]), .B(sum12[17][i12]), .Out(sum12[20][i12]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum12[18][i12]), .B(sum12[19][i12]), .Out(sum12[21][i12]));
      FP16_Add stage047(.A(sum12[20][i12]), .B(multi12[24][i12]), .Out(sum12[22][i12]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum12[21][i12]), .B(sum12[22][i12]), .Out(sum12[23][i12]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum12[23][i12]), .B(feature3Bias), .Out(data_11_array[j12][i12]));
    end
  endgenerate

  ////ROW 13
  generate
    localparam integer j13 = 13;
    for (i13 = 0; i13 < 24; i13 = i13 + 1)
    begin: addbit13
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j13+0][i13+0]), .Out(multi13[0][i13]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j13+0][i13+1]), .Out(multi13[1][i13]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j13+0][i13+2]), .Out(multi13[2][i13]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j13+0][i13+3]), .Out(multi13[3][i13]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j13+0][i13+4]), .Out(multi13[4][i13]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j13+1][i13+0]), .Out(multi13[5][i13]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j13+1][i13+1]), .Out(multi13[6][i13]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j13+1][i13+2]), .Out(multi13[7][i13]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j13+1][i13+3]), .Out(multi13[8][i13]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j13+1][i13+4]), .Out(multi13[9][i13]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j13+2][i13+0]), .Out(multi13[10][i13]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j13+2][i13+1]), .Out(multi13[11][i13]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j13+2][i13+2]), .Out(multi13[12][i13]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j13+2][i13+3]), .Out(multi13[13][i13]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j13+2][i13+4]), .Out(multi13[14][i13]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j13+3][i13+0]), .Out(multi13[15][i13]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j13+3][i13+1]), .Out(multi13[16][i13]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j13+3][i13+2]), .Out(multi13[17][i13]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j13+3][i13+3]), .Out(multi13[18][i13]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j13+3][i13+4]), .Out(multi13[19][i13]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j13+4][i13+0]), .Out(multi13[20][i13]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j13+4][i13+1]), .Out(multi13[21][i13]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j13+4][i13+2]), .Out(multi13[22][i13]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j13+4][i13+3]), .Out(multi13[23][i13]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j13+4][i13+4]), .Out(multi13[24][i13]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi13[0][i13]), .B(multi13[1][i13]), .Out(sum13[0][i13]));
      FP16_Add stage026(.A(multi13[2][i13]), .B(multi13[3][i13]), .Out(sum13[1][i13]));
      FP16_Add stage027(.A(multi13[4][i13]), .B(multi13[5][i13]), .Out(sum13[2][i13]));
      FP16_Add stage028(.A(multi13[6][i13]), .B(multi13[7][i13]), .Out(sum13[3][i13]));
      FP16_Add stage029(.A(multi13[8][i13]), .B(multi13[9][i13]), .Out(sum13[4][i13]));
      FP16_Add stage030(.A(multi13[10][i13]), .B(multi13[11][i13]), .Out(sum13[5][i13]));
      FP16_Add stage031(.A(multi13[12][i13]), .B(multi13[13][i13]), .Out(sum13[6][i13]));
      FP16_Add stage032(.A(multi13[14][i13]), .B(multi13[15][i13]), .Out(sum13[7][i13]));
      FP16_Add stage033(.A(multi13[16][i13]), .B(multi13[17][i13]), .Out(sum13[8][i13]));
      FP16_Add stage034(.A(multi13[18][i13]), .B(multi13[19][i13]), .Out(sum13[9][i13]));
      FP16_Add stage035(.A(multi13[20][i13]), .B(multi13[21][i13]), .Out(sum13[10][i13]));
      FP16_Add stage036(.A(multi13[22][i13]), .B(multi13[23][i13]), .Out(sum13[11][i13]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum13[0][i13]), .B(sum13[1][i13]), .Out(sum13[12][i13]));
      FP16_Add stage038(.A(sum13[2][i13]), .B(sum13[3][i13]), .Out(sum13[13][i13]));
      FP16_Add stage039(.A(sum13[4][i13]), .B(sum13[5][i13]), .Out(sum13[14][i13]));
      FP16_Add stage040(.A(sum13[6][i13]), .B(sum13[7][i13]), .Out(sum13[15][i13]));
      FP16_Add stage041(.A(sum13[8][i13]), .B(sum13[9][i13]), .Out(sum13[16][i13]));
      FP16_Add stage042(.A(sum13[10][i13]), .B(sum13[11][i13]), .Out(sum13[17][i13]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum13[12][i13]), .B(sum13[13][i13]), .Out(sum13[18][i13]));
      FP16_Add stage044(.A(sum13[14][i13]), .B(sum13[15][i13]), .Out(sum13[19][i13]));
      FP16_Add stage045(.A(sum13[16][i13]), .B(sum13[17][i13]), .Out(sum13[20][i13]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum13[18][i13]), .B(sum13[19][i13]), .Out(sum13[21][i13]));
      FP16_Add stage047(.A(sum13[20][i13]), .B(multi13[24][i13]), .Out(sum13[22][i13]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum13[21][i13]), .B(sum13[22][i13]), .Out(sum13[23][i13]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum13[23][i13]), .B(feature3Bias), .Out(data_11_array[j13][i13]));
    end
  endgenerate

  ////ROW 014
  generate
    localparam integer j14 = 14;
    for (i14 = 0; i14 < 24; i14 = i14 + 1)
    begin: addbit14
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j14+0][i14+0]), .Out(multi14[0][i14]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j14+0][i14+1]), .Out(multi14[1][i14]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j14+0][i14+2]), .Out(multi14[2][i14]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j14+0][i14+3]), .Out(multi14[3][i14]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j14+0][i14+4]), .Out(multi14[4][i14]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j14+1][i14+0]), .Out(multi14[5][i14]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j14+1][i14+1]), .Out(multi14[6][i14]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j14+1][i14+2]), .Out(multi14[7][i14]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j14+1][i14+3]), .Out(multi14[8][i14]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j14+1][i14+4]), .Out(multi14[9][i14]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j14+2][i14+0]), .Out(multi14[10][i14]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j14+2][i14+1]), .Out(multi14[11][i14]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j14+2][i14+2]), .Out(multi14[12][i14]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j14+2][i14+3]), .Out(multi14[13][i14]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j14+2][i14+4]), .Out(multi14[14][i14]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j14+3][i14+0]), .Out(multi14[15][i14]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j14+3][i14+1]), .Out(multi14[16][i14]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j14+3][i14+2]), .Out(multi14[17][i14]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j14+3][i14+3]), .Out(multi14[18][i14]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j14+3][i14+4]), .Out(multi14[19][i14]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j14+4][i14+0]), .Out(multi14[20][i14]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j14+4][i14+1]), .Out(multi14[21][i14]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j14+4][i14+2]), .Out(multi14[22][i14]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j14+4][i14+3]), .Out(multi14[23][i14]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j14+4][i14+4]), .Out(multi14[24][i14]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi14[0][i14]), .B(multi14[1][i14]), .Out(sum14[0][i14]));
      FP16_Add stage026(.A(multi14[2][i14]), .B(multi14[3][i14]), .Out(sum14[1][i14]));
      FP16_Add stage027(.A(multi14[4][i14]), .B(multi14[5][i14]), .Out(sum14[2][i14]));
      FP16_Add stage028(.A(multi14[6][i14]), .B(multi14[7][i14]), .Out(sum14[3][i14]));
      FP16_Add stage029(.A(multi14[8][i14]), .B(multi14[9][i14]), .Out(sum14[4][i14]));
      FP16_Add stage030(.A(multi14[10][i14]), .B(multi14[11][i14]), .Out(sum14[5][i14]));
      FP16_Add stage031(.A(multi14[12][i14]), .B(multi14[13][i14]), .Out(sum14[6][i14]));
      FP16_Add stage032(.A(multi14[14][i14]), .B(multi14[15][i14]), .Out(sum14[7][i14]));
      FP16_Add stage033(.A(multi14[16][i14]), .B(multi14[17][i14]), .Out(sum14[8][i14]));
      FP16_Add stage034(.A(multi14[18][i14]), .B(multi14[19][i14]), .Out(sum14[9][i14]));
      FP16_Add stage035(.A(multi14[20][i14]), .B(multi14[21][i14]), .Out(sum14[10][i14]));
      FP16_Add stage036(.A(multi14[22][i14]), .B(multi14[23][i14]), .Out(sum14[11][i14]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum14[0][i14]), .B(sum14[1][i14]), .Out(sum14[12][i14]));
      FP16_Add stage038(.A(sum14[2][i14]), .B(sum14[3][i14]), .Out(sum14[13][i14]));
      FP16_Add stage039(.A(sum14[4][i14]), .B(sum14[5][i14]), .Out(sum14[14][i14]));
      FP16_Add stage040(.A(sum14[6][i14]), .B(sum14[7][i14]), .Out(sum14[15][i14]));
      FP16_Add stage041(.A(sum14[8][i14]), .B(sum14[9][i14]), .Out(sum14[16][i14]));
      FP16_Add stage042(.A(sum14[10][i14]), .B(sum14[11][i14]), .Out(sum14[17][i14]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum14[12][i14]), .B(sum14[13][i14]), .Out(sum14[18][i14]));
      FP16_Add stage044(.A(sum14[14][i14]), .B(sum14[15][i14]), .Out(sum14[19][i14]));
      FP16_Add stage045(.A(sum14[16][i14]), .B(sum14[17][i14]), .Out(sum14[20][i14]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum14[18][i14]), .B(sum14[19][i14]), .Out(sum14[21][i14]));
      FP16_Add stage047(.A(sum14[20][i14]), .B(multi14[24][i14]), .Out(sum14[22][i14]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum14[21][i14]), .B(sum14[22][i14]), .Out(sum14[23][i14]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum14[23][i14]), .B(feature3Bias), .Out(data_11_array[j14][i14]));
    end
  endgenerate

  ////ROW 15
  generate
    localparam integer j15 = 15;
    for (i15 = 0; i15 < 24; i15 = i15 + 1)
    begin: addbit15
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j15+0][i15+0]), .Out(multi15[0][i15]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j15+0][i15+1]), .Out(multi15[1][i15]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j15+0][i15+2]), .Out(multi15[2][i15]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j15+0][i15+3]), .Out(multi15[3][i15]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j15+0][i15+4]), .Out(multi15[4][i15]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j15+1][i15+0]), .Out(multi15[5][i15]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j15+1][i15+1]), .Out(multi15[6][i15]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j15+1][i15+2]), .Out(multi15[7][i15]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j15+1][i15+3]), .Out(multi15[8][i15]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j15+1][i15+4]), .Out(multi15[9][i15]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j15+2][i15+0]), .Out(multi15[10][i15]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j15+2][i15+1]), .Out(multi15[11][i15]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j15+2][i15+2]), .Out(multi15[12][i15]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j15+2][i15+3]), .Out(multi15[13][i15]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j15+2][i15+4]), .Out(multi15[14][i15]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j15+3][i15+0]), .Out(multi15[15][i15]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j15+3][i15+1]), .Out(multi15[16][i15]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j15+3][i15+2]), .Out(multi15[17][i15]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j15+3][i15+3]), .Out(multi15[18][i15]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j15+3][i15+4]), .Out(multi15[19][i15]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j15+4][i15+0]), .Out(multi15[20][i15]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j15+4][i15+1]), .Out(multi15[21][i15]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j15+4][i15+2]), .Out(multi15[22][i15]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j15+4][i15+3]), .Out(multi15[23][i15]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j15+4][i15+4]), .Out(multi15[24][i15]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi15[0][i15]), .B(multi15[1][i15]), .Out(sum15[0][i15]));
      FP16_Add stage026(.A(multi15[2][i15]), .B(multi15[3][i15]), .Out(sum15[1][i15]));
      FP16_Add stage027(.A(multi15[4][i15]), .B(multi15[5][i15]), .Out(sum15[2][i15]));
      FP16_Add stage028(.A(multi15[6][i15]), .B(multi15[7][i15]), .Out(sum15[3][i15]));
      FP16_Add stage029(.A(multi15[8][i15]), .B(multi15[9][i15]), .Out(sum15[4][i15]));
      FP16_Add stage030(.A(multi15[10][i15]), .B(multi15[11][i15]), .Out(sum15[5][i15]));
      FP16_Add stage031(.A(multi15[12][i15]), .B(multi15[13][i15]), .Out(sum15[6][i15]));
      FP16_Add stage032(.A(multi15[14][i15]), .B(multi15[15][i15]), .Out(sum15[7][i15]));
      FP16_Add stage033(.A(multi15[16][i15]), .B(multi15[17][i15]), .Out(sum15[8][i15]));
      FP16_Add stage034(.A(multi15[18][i15]), .B(multi15[19][i15]), .Out(sum15[9][i15]));
      FP16_Add stage035(.A(multi15[20][i15]), .B(multi15[21][i15]), .Out(sum15[10][i15]));
      FP16_Add stage036(.A(multi15[22][i15]), .B(multi15[23][i15]), .Out(sum15[11][i15]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum15[0][i15]), .B(sum15[1][i15]), .Out(sum15[12][i15]));
      FP16_Add stage038(.A(sum15[2][i15]), .B(sum15[3][i15]), .Out(sum15[13][i15]));
      FP16_Add stage039(.A(sum15[4][i15]), .B(sum15[5][i15]), .Out(sum15[14][i15]));
      FP16_Add stage040(.A(sum15[6][i15]), .B(sum15[7][i15]), .Out(sum15[15][i15]));
      FP16_Add stage041(.A(sum15[8][i15]), .B(sum15[9][i15]), .Out(sum15[16][i15]));
      FP16_Add stage042(.A(sum15[10][i15]), .B(sum15[11][i15]), .Out(sum15[17][i15]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum15[12][i15]), .B(sum15[13][i15]), .Out(sum15[18][i15]));
      FP16_Add stage044(.A(sum15[14][i15]), .B(sum15[15][i15]), .Out(sum15[19][i15]));
      FP16_Add stage045(.A(sum15[16][i15]), .B(sum15[17][i15]), .Out(sum15[20][i15]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum15[18][i15]), .B(sum15[19][i15]), .Out(sum15[21][i15]));
      FP16_Add stage047(.A(sum15[20][i15]), .B(multi15[24][i15]), .Out(sum15[22][i15]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum15[21][i15]), .B(sum15[22][i15]), .Out(sum15[23][i15]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum15[23][i15]), .B(feature3Bias), .Out(data_11_array[j15][i15]));
    end
  endgenerate
  
  ////ROW 16
  generate
    localparam integer j16 = 16;
    for (i16 = 0; i16 < 24; i16 = i16 + 1)
    begin: addbit16
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j16+0][i16+0]), .Out(multi16[0][i16]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j16+0][i16+1]), .Out(multi16[1][i16]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j16+0][i16+2]), .Out(multi16[2][i16]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j16+0][i16+3]), .Out(multi16[3][i16]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j16+0][i16+4]), .Out(multi16[4][i16]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j16+1][i16+0]), .Out(multi16[5][i16]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j16+1][i16+1]), .Out(multi16[6][i16]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j16+1][i16+2]), .Out(multi16[7][i16]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j16+1][i16+3]), .Out(multi16[8][i16]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j16+1][i16+4]), .Out(multi16[9][i16]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j16+2][i16+0]), .Out(multi16[10][i16]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j16+2][i16+1]), .Out(multi16[11][i16]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j16+2][i16+2]), .Out(multi16[12][i16]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j16+2][i16+3]), .Out(multi16[13][i16]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j16+2][i16+4]), .Out(multi16[14][i16]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j16+3][i16+0]), .Out(multi16[15][i16]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j16+3][i16+1]), .Out(multi16[16][i16]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j16+3][i16+2]), .Out(multi16[17][i16]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j16+3][i16+3]), .Out(multi16[18][i16]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j16+3][i16+4]), .Out(multi16[19][i16]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j16+4][i16+0]), .Out(multi16[20][i16]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j16+4][i16+1]), .Out(multi16[21][i16]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j16+4][i16+2]), .Out(multi16[22][i16]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j16+4][i16+3]), .Out(multi16[23][i16]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j16+4][i16+4]), .Out(multi16[24][i16]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi16[0][i16]), .B(multi16[1][i16]), .Out(sum16[0][i16]));
      FP16_Add stage026(.A(multi16[2][i16]), .B(multi16[3][i16]), .Out(sum16[1][i16]));
      FP16_Add stage027(.A(multi16[4][i16]), .B(multi16[5][i16]), .Out(sum16[2][i16]));
      FP16_Add stage028(.A(multi16[6][i16]), .B(multi16[7][i16]), .Out(sum16[3][i16]));
      FP16_Add stage029(.A(multi16[8][i16]), .B(multi16[9][i16]), .Out(sum16[4][i16]));
      FP16_Add stage030(.A(multi16[10][i16]), .B(multi16[11][i16]), .Out(sum16[5][i16]));
      FP16_Add stage031(.A(multi16[12][i16]), .B(multi16[13][i16]), .Out(sum16[6][i16]));
      FP16_Add stage032(.A(multi16[14][i16]), .B(multi16[15][i16]), .Out(sum16[7][i16]));
      FP16_Add stage033(.A(multi16[16][i16]), .B(multi16[17][i16]), .Out(sum16[8][i16]));
      FP16_Add stage034(.A(multi16[18][i16]), .B(multi16[19][i16]), .Out(sum16[9][i16]));
      FP16_Add stage035(.A(multi16[20][i16]), .B(multi16[21][i16]), .Out(sum16[10][i16]));
      FP16_Add stage036(.A(multi16[22][i16]), .B(multi16[23][i16]), .Out(sum16[11][i16]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum16[0][i16]), .B(sum16[1][i16]), .Out(sum16[12][i16]));
      FP16_Add stage038(.A(sum16[2][i16]), .B(sum16[3][i16]), .Out(sum16[13][i16]));
      FP16_Add stage039(.A(sum16[4][i16]), .B(sum16[5][i16]), .Out(sum16[14][i16]));
      FP16_Add stage040(.A(sum16[6][i16]), .B(sum16[7][i16]), .Out(sum16[15][i16]));
      FP16_Add stage041(.A(sum16[8][i16]), .B(sum16[9][i16]), .Out(sum16[16][i16]));
      FP16_Add stage042(.A(sum16[10][i16]), .B(sum16[11][i16]), .Out(sum16[17][i16]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum16[12][i16]), .B(sum16[13][i16]), .Out(sum16[18][i16]));
      FP16_Add stage044(.A(sum16[14][i16]), .B(sum16[15][i16]), .Out(sum16[19][i16]));
      FP16_Add stage045(.A(sum16[16][i16]), .B(sum16[17][i16]), .Out(sum16[20][i16]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum16[18][i16]), .B(sum16[19][i16]), .Out(sum16[21][i16]));
      FP16_Add stage047(.A(sum16[20][i16]), .B(multi16[24][i16]), .Out(sum16[22][i16]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum16[21][i16]), .B(sum16[22][i16]), .Out(sum16[23][i16]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum16[23][i16]), .B(feature3Bias), .Out(data_11_array[j16][i16]));
    end
  endgenerate
  
  ////ROW 17
  generate
    localparam integer j17 = 17;
    for (i17 = 0; i17 < 24; i17 = i17 + 1)
    begin: addbit17
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j17+0][i17+0]), .Out(multi17[0][i17]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j17+0][i17+1]), .Out(multi17[1][i17]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j17+0][i17+2]), .Out(multi17[2][i17]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j17+0][i17+3]), .Out(multi17[3][i17]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j17+0][i17+4]), .Out(multi17[4][i17]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j17+1][i17+0]), .Out(multi17[5][i17]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j17+1][i17+1]), .Out(multi17[6][i17]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j17+1][i17+2]), .Out(multi17[7][i17]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j17+1][i17+3]), .Out(multi17[8][i17]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j17+1][i17+4]), .Out(multi17[9][i17]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j17+2][i17+0]), .Out(multi17[10][i17]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j17+2][i17+1]), .Out(multi17[11][i17]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j17+2][i17+2]), .Out(multi17[12][i17]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j17+2][i17+3]), .Out(multi17[13][i17]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j17+2][i17+4]), .Out(multi17[14][i17]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j17+3][i17+0]), .Out(multi17[15][i17]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j17+3][i17+1]), .Out(multi17[16][i17]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j17+3][i17+2]), .Out(multi17[17][i17]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j17+3][i17+3]), .Out(multi17[18][i17]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j17+3][i17+4]), .Out(multi17[19][i17]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j17+4][i17+0]), .Out(multi17[20][i17]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j17+4][i17+1]), .Out(multi17[21][i17]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j17+4][i17+2]), .Out(multi17[22][i17]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j17+4][i17+3]), .Out(multi17[23][i17]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j17+4][i17+4]), .Out(multi17[24][i17]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi17[0][i17]), .B(multi17[1][i17]), .Out(sum17[0][i17]));
      FP16_Add stage026(.A(multi17[2][i17]), .B(multi17[3][i17]), .Out(sum17[1][i17]));
      FP16_Add stage027(.A(multi17[4][i17]), .B(multi17[5][i17]), .Out(sum17[2][i17]));
      FP16_Add stage028(.A(multi17[6][i17]), .B(multi17[7][i17]), .Out(sum17[3][i17]));
      FP16_Add stage029(.A(multi17[8][i17]), .B(multi17[9][i17]), .Out(sum17[4][i17]));
      FP16_Add stage030(.A(multi17[10][i17]), .B(multi17[11][i17]), .Out(sum17[5][i17]));
      FP16_Add stage031(.A(multi17[12][i17]), .B(multi17[13][i17]), .Out(sum17[6][i17]));
      FP16_Add stage032(.A(multi17[14][i17]), .B(multi17[15][i17]), .Out(sum17[7][i17]));
      FP16_Add stage033(.A(multi17[16][i17]), .B(multi17[17][i17]), .Out(sum17[8][i17]));
      FP16_Add stage034(.A(multi17[18][i17]), .B(multi17[19][i17]), .Out(sum17[9][i17]));
      FP16_Add stage035(.A(multi17[20][i17]), .B(multi17[21][i17]), .Out(sum17[10][i17]));
      FP16_Add stage036(.A(multi17[22][i17]), .B(multi17[23][i17]), .Out(sum17[11][i17]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum17[0][i17]), .B(sum17[1][i17]), .Out(sum17[12][i17]));
      FP16_Add stage038(.A(sum17[2][i17]), .B(sum17[3][i17]), .Out(sum17[13][i17]));
      FP16_Add stage039(.A(sum17[4][i17]), .B(sum17[5][i17]), .Out(sum17[14][i17]));
      FP16_Add stage040(.A(sum17[6][i17]), .B(sum17[7][i17]), .Out(sum17[15][i17]));
      FP16_Add stage041(.A(sum17[8][i17]), .B(sum17[9][i17]), .Out(sum17[16][i17]));
      FP16_Add stage042(.A(sum17[10][i17]), .B(sum17[11][i17]), .Out(sum17[17][i17]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum17[12][i17]), .B(sum17[13][i17]), .Out(sum17[18][i17]));
      FP16_Add stage044(.A(sum17[14][i17]), .B(sum17[15][i17]), .Out(sum17[19][i17]));
      FP16_Add stage045(.A(sum17[16][i17]), .B(sum17[17][i17]), .Out(sum17[20][i17]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum17[18][i17]), .B(sum17[19][i17]), .Out(sum17[21][i17]));
      FP16_Add stage047(.A(sum17[20][i17]), .B(multi17[24][i17]), .Out(sum17[22][i17]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum17[21][i17]), .B(sum17[22][i17]), .Out(sum17[23][i17]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum17[23][i17]), .B(feature3Bias), .Out(data_11_array[j17][i17]));
    end
  endgenerate

////ROW 18
  generate
    localparam integer j18 = 18;
    for (i18 = 0; i18 < 24; i18 = i18 + 1)
    begin: addbit18
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j18+0][i18+0]), .Out(multi18[0][i18]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j18+0][i18+1]), .Out(multi18[1][i18]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j18+0][i18+2]), .Out(multi18[2][i18]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j18+0][i18+3]), .Out(multi18[3][i18]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j18+0][i18+4]), .Out(multi18[4][i18]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j18+1][i18+0]), .Out(multi18[5][i18]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j18+1][i18+1]), .Out(multi18[6][i18]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j18+1][i18+2]), .Out(multi18[7][i18]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j18+1][i18+3]), .Out(multi18[8][i18]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j18+1][i18+4]), .Out(multi18[9][i18]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j18+2][i18+0]), .Out(multi18[10][i18]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j18+2][i18+1]), .Out(multi18[11][i18]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j18+2][i18+2]), .Out(multi18[12][i18]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j18+2][i18+3]), .Out(multi18[13][i18]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j18+2][i18+4]), .Out(multi18[14][i18]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j18+3][i18+0]), .Out(multi18[15][i18]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j18+3][i18+1]), .Out(multi18[16][i18]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j18+3][i18+2]), .Out(multi18[17][i18]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j18+3][i18+3]), .Out(multi18[18][i18]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j18+3][i18+4]), .Out(multi18[19][i18]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j18+4][i18+0]), .Out(multi18[20][i18]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j18+4][i18+1]), .Out(multi18[21][i18]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j18+4][i18+2]), .Out(multi18[22][i18]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j18+4][i18+3]), .Out(multi18[23][i18]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j18+4][i18+4]), .Out(multi18[24][i18]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi18[0][i18]), .B(multi18[1][i18]), .Out(sum18[0][i18]));
      FP16_Add stage026(.A(multi18[2][i18]), .B(multi18[3][i18]), .Out(sum18[1][i18]));
      FP16_Add stage027(.A(multi18[4][i18]), .B(multi18[5][i18]), .Out(sum18[2][i18]));
      FP16_Add stage028(.A(multi18[6][i18]), .B(multi18[7][i18]), .Out(sum18[3][i18]));
      FP16_Add stage029(.A(multi18[8][i18]), .B(multi18[9][i18]), .Out(sum18[4][i18]));
      FP16_Add stage030(.A(multi18[10][i18]), .B(multi18[11][i18]), .Out(sum18[5][i18]));
      FP16_Add stage031(.A(multi18[12][i18]), .B(multi18[13][i18]), .Out(sum18[6][i18]));
      FP16_Add stage032(.A(multi18[14][i18]), .B(multi18[15][i18]), .Out(sum18[7][i18]));
      FP16_Add stage033(.A(multi18[16][i18]), .B(multi18[17][i18]), .Out(sum18[8][i18]));
      FP16_Add stage034(.A(multi18[18][i18]), .B(multi18[19][i18]), .Out(sum18[9][i18]));
      FP16_Add stage035(.A(multi18[20][i18]), .B(multi18[21][i18]), .Out(sum18[10][i18]));
      FP16_Add stage036(.A(multi18[22][i18]), .B(multi18[23][i18]), .Out(sum18[11][i18]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum18[0][i18]), .B(sum18[1][i18]), .Out(sum18[12][i18]));
      FP16_Add stage038(.A(sum18[2][i18]), .B(sum18[3][i18]), .Out(sum18[13][i18]));
      FP16_Add stage039(.A(sum18[4][i18]), .B(sum18[5][i18]), .Out(sum18[14][i18]));
      FP16_Add stage040(.A(sum18[6][i18]), .B(sum18[7][i18]), .Out(sum18[15][i18]));
      FP16_Add stage041(.A(sum18[8][i18]), .B(sum18[9][i18]), .Out(sum18[16][i18]));
      FP16_Add stage042(.A(sum18[10][i18]), .B(sum18[11][i18]), .Out(sum18[17][i18]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum18[12][i18]), .B(sum18[13][i18]), .Out(sum18[18][i18]));
      FP16_Add stage044(.A(sum18[14][i18]), .B(sum18[15][i18]), .Out(sum18[19][i18]));
      FP16_Add stage045(.A(sum18[16][i18]), .B(sum18[17][i18]), .Out(sum18[20][i18]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum18[18][i18]), .B(sum18[19][i18]), .Out(sum18[21][i18]));
      FP16_Add stage047(.A(sum18[20][i18]), .B(multi18[24][i18]), .Out(sum18[22][i18]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum18[21][i18]), .B(sum18[22][i18]), .Out(sum18[23][i18]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum18[23][i18]), .B(feature3Bias), .Out(data_11_array[j18][i18]));
    end
  endgenerate

////ROW 19
  generate
    localparam integer j19 = 19;
    for (i19 = 0; i19 < 24; i19 = i19 + 1)
    begin: addbit19
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j19+0][i19+0]), .Out(multi19[0][i19]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j19+0][i19+1]), .Out(multi19[1][i19]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j19+0][i19+2]), .Out(multi19[2][i19]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j19+0][i19+3]), .Out(multi19[3][i19]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j19+0][i19+4]), .Out(multi19[4][i19]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j19+1][i19+0]), .Out(multi19[5][i19]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j19+1][i19+1]), .Out(multi19[6][i19]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j19+1][i19+2]), .Out(multi19[7][i19]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j19+1][i19+3]), .Out(multi19[8][i19]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j19+1][i19+4]), .Out(multi19[9][i19]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j19+2][i19+0]), .Out(multi19[10][i19]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j19+2][i19+1]), .Out(multi19[11][i19]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j19+2][i19+2]), .Out(multi19[12][i19]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j19+2][i19+3]), .Out(multi19[13][i19]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j19+2][i19+4]), .Out(multi19[14][i19]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j19+3][i19+0]), .Out(multi19[15][i19]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j19+3][i19+1]), .Out(multi19[16][i19]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j19+3][i19+2]), .Out(multi19[17][i19]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j19+3][i19+3]), .Out(multi19[18][i19]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j19+3][i19+4]), .Out(multi19[19][i19]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j19+4][i19+0]), .Out(multi19[20][i19]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j19+4][i19+1]), .Out(multi19[21][i19]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j19+4][i19+2]), .Out(multi19[22][i19]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j19+4][i19+3]), .Out(multi19[23][i19]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j19+4][i19+4]), .Out(multi19[24][i19]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi19[0][i19]), .B(multi19[1][i19]), .Out(sum19[0][i19]));
      FP16_Add stage026(.A(multi19[2][i19]), .B(multi19[3][i19]), .Out(sum19[1][i19]));
      FP16_Add stage027(.A(multi19[4][i19]), .B(multi19[5][i19]), .Out(sum19[2][i19]));
      FP16_Add stage028(.A(multi19[6][i19]), .B(multi19[7][i19]), .Out(sum19[3][i19]));
      FP16_Add stage029(.A(multi19[8][i19]), .B(multi19[9][i19]), .Out(sum19[4][i19]));
      FP16_Add stage030(.A(multi19[10][i19]), .B(multi19[11][i19]), .Out(sum19[5][i19]));
      FP16_Add stage031(.A(multi19[12][i19]), .B(multi19[13][i19]), .Out(sum19[6][i19]));
      FP16_Add stage032(.A(multi19[14][i19]), .B(multi19[15][i19]), .Out(sum19[7][i19]));
      FP16_Add stage033(.A(multi19[16][i19]), .B(multi19[17][i19]), .Out(sum19[8][i19]));
      FP16_Add stage034(.A(multi19[18][i19]), .B(multi19[19][i19]), .Out(sum19[9][i19]));
      FP16_Add stage035(.A(multi19[20][i19]), .B(multi19[21][i19]), .Out(sum19[10][i19]));
      FP16_Add stage036(.A(multi19[22][i19]), .B(multi19[23][i19]), .Out(sum19[11][i19]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum19[0][i19]), .B(sum19[1][i19]), .Out(sum19[12][i19]));
      FP16_Add stage038(.A(sum19[2][i19]), .B(sum19[3][i19]), .Out(sum19[13][i19]));
      FP16_Add stage039(.A(sum19[4][i19]), .B(sum19[5][i19]), .Out(sum19[14][i19]));
      FP16_Add stage040(.A(sum19[6][i19]), .B(sum19[7][i19]), .Out(sum19[15][i19]));
      FP16_Add stage041(.A(sum19[8][i19]), .B(sum19[9][i19]), .Out(sum19[16][i19]));
      FP16_Add stage042(.A(sum19[10][i19]), .B(sum19[11][i19]), .Out(sum19[17][i19]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum19[12][i19]), .B(sum19[13][i19]), .Out(sum19[18][i19]));
      FP16_Add stage044(.A(sum19[14][i19]), .B(sum19[15][i19]), .Out(sum19[19][i19]));
      FP16_Add stage045(.A(sum19[16][i19]), .B(sum19[17][i19]), .Out(sum19[20][i19]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum19[18][i19]), .B(sum19[19][i19]), .Out(sum19[21][i19]));
      FP16_Add stage047(.A(sum19[20][i19]), .B(multi19[24][i19]), .Out(sum19[22][i19]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum19[21][i19]), .B(sum19[22][i19]), .Out(sum19[23][i19]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum19[23][i19]), .B(feature3Bias), .Out(data_11_array[j19][i19]));
    end
  endgenerate

////ROW 20
  generate
    localparam integer j20 = 20;
    for (i20 = 0; i20 < 24; i20 = i20 + 1)
    begin: addbit20
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j20+0][i20+0]), .Out(multi20[0][i20]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j20+0][i20+1]), .Out(multi20[1][i20]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j20+0][i20+2]), .Out(multi20[2][i20]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j20+0][i20+3]), .Out(multi20[3][i20]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j20+0][i20+4]), .Out(multi20[4][i20]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j20+1][i20+0]), .Out(multi20[5][i20]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j20+1][i20+1]), .Out(multi20[6][i20]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j20+1][i20+2]), .Out(multi20[7][i20]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j20+1][i20+3]), .Out(multi20[8][i20]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j20+1][i20+4]), .Out(multi20[9][i20]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j20+2][i20+0]), .Out(multi20[10][i20]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j20+2][i20+1]), .Out(multi20[11][i20]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j20+2][i20+2]), .Out(multi20[12][i20]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j20+2][i20+3]), .Out(multi20[13][i20]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j20+2][i20+4]), .Out(multi20[14][i20]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j20+3][i20+0]), .Out(multi20[15][i20]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j20+3][i20+1]), .Out(multi20[16][i20]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j20+3][i20+2]), .Out(multi20[17][i20]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j20+3][i20+3]), .Out(multi20[18][i20]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j20+3][i20+4]), .Out(multi20[19][i20]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j20+4][i20+0]), .Out(multi20[20][i20]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j20+4][i20+1]), .Out(multi20[21][i20]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j20+4][i20+2]), .Out(multi20[22][i20]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j20+4][i20+3]), .Out(multi20[23][i20]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j20+4][i20+4]), .Out(multi20[24][i20]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi20[0][i20]), .B(multi20[1][i20]), .Out(sum20[0][i20]));
      FP16_Add stage026(.A(multi20[2][i20]), .B(multi20[3][i20]), .Out(sum20[1][i20]));
      FP16_Add stage027(.A(multi20[4][i20]), .B(multi20[5][i20]), .Out(sum20[2][i20]));
      FP16_Add stage028(.A(multi20[6][i20]), .B(multi20[7][i20]), .Out(sum20[3][i20]));
      FP16_Add stage029(.A(multi20[8][i20]), .B(multi20[9][i20]), .Out(sum20[4][i20]));
      FP16_Add stage030(.A(multi20[10][i20]), .B(multi20[11][i20]), .Out(sum20[5][i20]));
      FP16_Add stage031(.A(multi20[12][i20]), .B(multi20[13][i20]), .Out(sum20[6][i20]));
      FP16_Add stage032(.A(multi20[14][i20]), .B(multi20[15][i20]), .Out(sum20[7][i20]));
      FP16_Add stage033(.A(multi20[16][i20]), .B(multi20[17][i20]), .Out(sum20[8][i20]));
      FP16_Add stage034(.A(multi20[18][i20]), .B(multi20[19][i20]), .Out(sum20[9][i20]));
      FP16_Add stage035(.A(multi20[20][i20]), .B(multi20[21][i20]), .Out(sum20[10][i20]));
      FP16_Add stage036(.A(multi20[22][i20]), .B(multi20[23][i20]), .Out(sum20[11][i20]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum20[0][i20]), .B(sum20[1][i20]), .Out(sum20[12][i20]));
      FP16_Add stage038(.A(sum20[2][i20]), .B(sum20[3][i20]), .Out(sum20[13][i20]));
      FP16_Add stage039(.A(sum20[4][i20]), .B(sum20[5][i20]), .Out(sum20[14][i20]));
      FP16_Add stage040(.A(sum20[6][i20]), .B(sum20[7][i20]), .Out(sum20[15][i20]));
      FP16_Add stage041(.A(sum20[8][i20]), .B(sum20[9][i20]), .Out(sum20[16][i20]));
      FP16_Add stage042(.A(sum20[10][i20]), .B(sum20[11][i20]), .Out(sum20[17][i20]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum20[12][i20]), .B(sum20[13][i20]), .Out(sum20[18][i20]));
      FP16_Add stage044(.A(sum20[14][i20]), .B(sum20[15][i20]), .Out(sum20[19][i20]));
      FP16_Add stage045(.A(sum20[16][i20]), .B(sum20[17][i20]), .Out(sum20[20][i20]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum20[18][i20]), .B(sum20[19][i20]), .Out(sum20[21][i20]));
      FP16_Add stage047(.A(sum20[20][i20]), .B(multi20[24][i20]), .Out(sum20[22][i20]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum20[21][i20]), .B(sum20[22][i20]), .Out(sum20[23][i20]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum20[23][i20]), .B(feature3Bias), .Out(data_11_array[j20][i20]));
    end
  endgenerate

////ROW 21
  generate
    localparam integer j21 = 21;
    for (i21 = 0; i21 < 24; i21 = i21 + 1)
    begin: addbit21
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j21+0][i21+0]), .Out(multi21[0][i21]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j21+0][i21+1]), .Out(multi21[1][i21]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j21+0][i21+2]), .Out(multi21[2][i21]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j21+0][i21+3]), .Out(multi21[3][i21]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j21+0][i21+4]), .Out(multi21[4][i21]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j21+1][i21+0]), .Out(multi21[5][i21]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j21+1][i21+1]), .Out(multi21[6][i21]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j21+1][i21+2]), .Out(multi21[7][i21]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j21+1][i21+3]), .Out(multi21[8][i21]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j21+1][i21+4]), .Out(multi21[9][i21]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j21+2][i21+0]), .Out(multi21[10][i21]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j21+2][i21+1]), .Out(multi21[11][i21]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j21+2][i21+2]), .Out(multi21[12][i21]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j21+2][i21+3]), .Out(multi21[13][i21]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j21+2][i21+4]), .Out(multi21[14][i21]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j21+3][i21+0]), .Out(multi21[15][i21]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j21+3][i21+1]), .Out(multi21[16][i21]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j21+3][i21+2]), .Out(multi21[17][i21]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j21+3][i21+3]), .Out(multi21[18][i21]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j21+3][i21+4]), .Out(multi21[19][i21]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j21+4][i21+0]), .Out(multi21[20][i21]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j21+4][i21+1]), .Out(multi21[21][i21]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j21+4][i21+2]), .Out(multi21[22][i21]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j21+4][i21+3]), .Out(multi21[23][i21]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j21+4][i21+4]), .Out(multi21[24][i21]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi21[0][i21]), .B(multi21[1][i21]), .Out(sum21[0][i21]));
      FP16_Add stage026(.A(multi21[2][i21]), .B(multi21[3][i21]), .Out(sum21[1][i21]));
      FP16_Add stage027(.A(multi21[4][i21]), .B(multi21[5][i21]), .Out(sum21[2][i21]));
      FP16_Add stage028(.A(multi21[6][i21]), .B(multi21[7][i21]), .Out(sum21[3][i21]));
      FP16_Add stage029(.A(multi21[8][i21]), .B(multi21[9][i21]), .Out(sum21[4][i21]));
      FP16_Add stage030(.A(multi21[10][i21]), .B(multi21[11][i21]), .Out(sum21[5][i21]));
      FP16_Add stage031(.A(multi21[12][i21]), .B(multi21[13][i21]), .Out(sum21[6][i21]));
      FP16_Add stage032(.A(multi21[14][i21]), .B(multi21[15][i21]), .Out(sum21[7][i21]));
      FP16_Add stage033(.A(multi21[16][i21]), .B(multi21[17][i21]), .Out(sum21[8][i21]));
      FP16_Add stage034(.A(multi21[18][i21]), .B(multi21[19][i21]), .Out(sum21[9][i21]));
      FP16_Add stage035(.A(multi21[20][i21]), .B(multi21[21][i21]), .Out(sum21[10][i21]));
      FP16_Add stage036(.A(multi21[22][i21]), .B(multi21[23][i21]), .Out(sum21[11][i21]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum21[0][i21]), .B(sum21[1][i21]), .Out(sum21[12][i21]));
      FP16_Add stage038(.A(sum21[2][i21]), .B(sum21[3][i21]), .Out(sum21[13][i21]));
      FP16_Add stage039(.A(sum21[4][i21]), .B(sum21[5][i21]), .Out(sum21[14][i21]));
      FP16_Add stage040(.A(sum21[6][i21]), .B(sum21[7][i21]), .Out(sum21[15][i21]));
      FP16_Add stage041(.A(sum21[8][i21]), .B(sum21[9][i21]), .Out(sum21[16][i21]));
      FP16_Add stage042(.A(sum21[10][i21]), .B(sum21[11][i21]), .Out(sum21[17][i21]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum21[12][i21]), .B(sum21[13][i21]), .Out(sum21[18][i21]));
      FP16_Add stage044(.A(sum21[14][i21]), .B(sum21[15][i21]), .Out(sum21[19][i21]));
      FP16_Add stage045(.A(sum21[16][i21]), .B(sum21[17][i21]), .Out(sum21[20][i21]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum21[18][i21]), .B(sum21[19][i21]), .Out(sum21[21][i21]));
      FP16_Add stage047(.A(sum21[20][i21]), .B(multi21[24][i21]), .Out(sum21[22][i21]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum21[21][i21]), .B(sum21[22][i21]), .Out(sum21[23][i21]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum21[23][i21]), .B(feature3Bias), .Out(data_11_array[j21][i21]));
    end
  endgenerate

////ROW 22
  generate
    localparam integer j22 = 22;
    for (i22 = 0; i22 < 24; i22 = i22 + 1)
    begin: addbit22
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j22+0][i22+0]), .Out(multi22[0][i22]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j22+0][i22+1]), .Out(multi22[1][i22]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j22+0][i22+2]), .Out(multi22[2][i22]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j22+0][i22+3]), .Out(multi22[3][i22]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j22+0][i22+4]), .Out(multi22[4][i22]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j22+1][i22+0]), .Out(multi22[5][i22]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j22+1][i22+1]), .Out(multi22[6][i22]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j22+1][i22+2]), .Out(multi22[7][i22]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j22+1][i22+3]), .Out(multi22[8][i22]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j22+1][i22+4]), .Out(multi22[9][i22]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j22+2][i22+0]), .Out(multi22[10][i22]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j22+2][i22+1]), .Out(multi22[11][i22]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j22+2][i22+2]), .Out(multi22[12][i22]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j22+2][i22+3]), .Out(multi22[13][i22]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j22+2][i22+4]), .Out(multi22[14][i22]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j22+3][i22+0]), .Out(multi22[15][i22]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j22+3][i22+1]), .Out(multi22[16][i22]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j22+3][i22+2]), .Out(multi22[17][i22]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j22+3][i22+3]), .Out(multi22[18][i22]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j22+3][i22+4]), .Out(multi22[19][i22]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j22+4][i22+0]), .Out(multi22[20][i22]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j22+4][i22+1]), .Out(multi22[21][i22]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j22+4][i22+2]), .Out(multi22[22][i22]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j22+4][i22+3]), .Out(multi22[23][i22]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j22+4][i22+4]), .Out(multi22[24][i22]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi22[0][i22]), .B(multi22[1][i22]), .Out(sum22[0][i22]));
      FP16_Add stage026(.A(multi22[2][i22]), .B(multi22[3][i22]), .Out(sum22[1][i22]));
      FP16_Add stage027(.A(multi22[4][i22]), .B(multi22[5][i22]), .Out(sum22[2][i22]));
      FP16_Add stage028(.A(multi22[6][i22]), .B(multi22[7][i22]), .Out(sum22[3][i22]));
      FP16_Add stage029(.A(multi22[8][i22]), .B(multi22[9][i22]), .Out(sum22[4][i22]));
      FP16_Add stage030(.A(multi22[10][i22]), .B(multi22[11][i22]), .Out(sum22[5][i22]));
      FP16_Add stage031(.A(multi22[12][i22]), .B(multi22[13][i22]), .Out(sum22[6][i22]));
      FP16_Add stage032(.A(multi22[14][i22]), .B(multi22[15][i22]), .Out(sum22[7][i22]));
      FP16_Add stage033(.A(multi22[16][i22]), .B(multi22[17][i22]), .Out(sum22[8][i22]));
      FP16_Add stage034(.A(multi22[18][i22]), .B(multi22[19][i22]), .Out(sum22[9][i22]));
      FP16_Add stage035(.A(multi22[20][i22]), .B(multi22[21][i22]), .Out(sum22[10][i22]));
      FP16_Add stage036(.A(multi22[22][i22]), .B(multi22[23][i22]), .Out(sum22[11][i22]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum22[0][i22]), .B(sum22[1][i22]), .Out(sum22[12][i22]));
      FP16_Add stage038(.A(sum22[2][i22]), .B(sum22[3][i22]), .Out(sum22[13][i22]));
      FP16_Add stage039(.A(sum22[4][i22]), .B(sum22[5][i22]), .Out(sum22[14][i22]));
      FP16_Add stage040(.A(sum22[6][i22]), .B(sum22[7][i22]), .Out(sum22[15][i22]));
      FP16_Add stage041(.A(sum22[8][i22]), .B(sum22[9][i22]), .Out(sum22[16][i22]));
      FP16_Add stage042(.A(sum22[10][i22]), .B(sum22[11][i22]), .Out(sum22[17][i22]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum22[12][i22]), .B(sum22[13][i22]), .Out(sum22[18][i22]));
      FP16_Add stage044(.A(sum22[14][i22]), .B(sum22[15][i22]), .Out(sum22[19][i22]));
      FP16_Add stage045(.A(sum22[16][i22]), .B(sum22[17][i22]), .Out(sum22[20][i22]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum22[18][i22]), .B(sum22[19][i22]), .Out(sum22[21][i22]));
      FP16_Add stage047(.A(sum22[20][i22]), .B(multi22[24][i22]), .Out(sum22[22][i22]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum22[21][i22]), .B(sum22[22][i22]), .Out(sum22[23][i22]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum22[23][i22]), .B(feature3Bias), .Out(data_11_array[j22][i22]));
    end
  endgenerate

////ROW 23
  generate
    localparam integer j23 = 23;
    for (i23 = 0; i23 < 24; i23 = i23 + 1)
    begin: addbit23
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature3Weight_0), .B(data_array[j23+0][i23+0]), .Out(multi23[0][i23]));
      FP16_Multiply stage01(.A(feature3Weight_1), .B(data_array[j23+0][i23+1]), .Out(multi23[1][i23]));
      FP16_Multiply stage02(.A(feature3Weight_2), .B(data_array[j23+0][i23+2]), .Out(multi23[2][i23]));
      FP16_Multiply stage03(.A(feature3Weight_3), .B(data_array[j23+0][i23+3]), .Out(multi23[3][i23]));
      FP16_Multiply stage04(.A(feature3Weight_4), .B(data_array[j23+0][i23+4]), .Out(multi23[4][i23]));
      FP16_Multiply stage05(.A(feature3Weight_5), .B(data_array[j23+1][i23+0]), .Out(multi23[5][i23]));
      FP16_Multiply stage06(.A(feature3Weight_6), .B(data_array[j23+1][i23+1]), .Out(multi23[6][i23]));
      FP16_Multiply stage07(.A(feature3Weight_7), .B(data_array[j23+1][i23+2]), .Out(multi23[7][i23]));
      FP16_Multiply stage08(.A(feature3Weight_8), .B(data_array[j23+1][i23+3]), .Out(multi23[8][i23]));
      FP16_Multiply stage09(.A(feature3Weight_9), .B(data_array[j23+1][i23+4]), .Out(multi23[9][i23]));
      FP16_Multiply stage010(.A(feature3Weight_10), .B(data_array[j23+2][i23+0]), .Out(multi23[10][i23]));
      FP16_Multiply stage011(.A(feature3Weight_11), .B(data_array[j23+2][i23+1]), .Out(multi23[11][i23]));
      FP16_Multiply stage012(.A(feature3Weight_12), .B(data_array[j23+2][i23+2]), .Out(multi23[12][i23]));
      FP16_Multiply stage013(.A(feature3Weight_13), .B(data_array[j23+2][i23+3]), .Out(multi23[13][i23]));
      FP16_Multiply stage014(.A(feature3Weight_14), .B(data_array[j23+2][i23+4]), .Out(multi23[14][i23]));
      FP16_Multiply stage015(.A(feature3Weight_15), .B(data_array[j23+3][i23+0]), .Out(multi23[15][i23]));
      FP16_Multiply stage016(.A(feature3Weight_16), .B(data_array[j23+3][i23+1]), .Out(multi23[16][i23]));
      FP16_Multiply stage017(.A(feature3Weight_17), .B(data_array[j23+3][i23+2]), .Out(multi23[17][i23]));
      FP16_Multiply stage018(.A(feature3Weight_18), .B(data_array[j23+3][i23+3]), .Out(multi23[18][i23]));
      FP16_Multiply stage019(.A(feature3Weight_19), .B(data_array[j23+3][i23+4]), .Out(multi23[19][i23]));
      FP16_Multiply stage020(.A(feature3Weight_20), .B(data_array[j23+4][i23+0]), .Out(multi23[20][i23]));
      FP16_Multiply stage021(.A(feature3Weight_21), .B(data_array[j23+4][i23+1]), .Out(multi23[21][i23]));
      FP16_Multiply stage022(.A(feature3Weight_22), .B(data_array[j23+4][i23+2]), .Out(multi23[22][i23]));
      FP16_Multiply stage023(.A(feature3Weight_23), .B(data_array[j23+4][i23+3]), .Out(multi23[23][i23]));
      FP16_Multiply stage024(.A(feature3Weight_24), .B(data_array[j23+4][i23+4]), .Out(multi23[24][i23]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi23[0][i23]), .B(multi23[1][i23]), .Out(sum23[0][i23]));
      FP16_Add stage026(.A(multi23[2][i23]), .B(multi23[3][i23]), .Out(sum23[1][i23]));
      FP16_Add stage027(.A(multi23[4][i23]), .B(multi23[5][i23]), .Out(sum23[2][i23]));
      FP16_Add stage028(.A(multi23[6][i23]), .B(multi23[7][i23]), .Out(sum23[3][i23]));
      FP16_Add stage029(.A(multi23[8][i23]), .B(multi23[9][i23]), .Out(sum23[4][i23]));
      FP16_Add stage030(.A(multi23[10][i23]), .B(multi23[11][i23]), .Out(sum23[5][i23]));
      FP16_Add stage031(.A(multi23[12][i23]), .B(multi23[13][i23]), .Out(sum23[6][i23]));
      FP16_Add stage032(.A(multi23[14][i23]), .B(multi23[15][i23]), .Out(sum23[7][i23]));
      FP16_Add stage033(.A(multi23[16][i23]), .B(multi23[17][i23]), .Out(sum23[8][i23]));
      FP16_Add stage034(.A(multi23[18][i23]), .B(multi23[19][i23]), .Out(sum23[9][i23]));
      FP16_Add stage035(.A(multi23[20][i23]), .B(multi23[21][i23]), .Out(sum23[10][i23]));
      FP16_Add stage036(.A(multi23[22][i23]), .B(multi23[23][i23]), .Out(sum23[11][i23]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum23[0][i23]), .B(sum23[1][i23]), .Out(sum23[12][i23]));
      FP16_Add stage038(.A(sum23[2][i23]), .B(sum23[3][i23]), .Out(sum23[13][i23]));
      FP16_Add stage039(.A(sum23[4][i23]), .B(sum23[5][i23]), .Out(sum23[14][i23]));
      FP16_Add stage040(.A(sum23[6][i23]), .B(sum23[7][i23]), .Out(sum23[15][i23]));
      FP16_Add stage041(.A(sum23[8][i23]), .B(sum23[9][i23]), .Out(sum23[16][i23]));
      FP16_Add stage042(.A(sum23[10][i23]), .B(sum23[11][i23]), .Out(sum23[17][i23]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum23[12][i23]), .B(sum23[13][i23]), .Out(sum23[18][i23]));
      FP16_Add stage044(.A(sum23[14][i23]), .B(sum23[15][i23]), .Out(sum23[19][i23]));
      FP16_Add stage045(.A(sum23[16][i23]), .B(sum23[17][i23]), .Out(sum23[20][i23]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum23[18][i23]), .B(sum23[19][i23]), .Out(sum23[21][i23]));
      FP16_Add stage047(.A(sum23[20][i23]), .B(multi23[24][i23]), .Out(sum23[22][i23]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum23[21][i23]), .B(sum23[22][i23]), .Out(sum23[23][i23]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum23[23][i23]), .B(feature3Bias), .Out(data_11_array[j23][i23]));
    end
  endgenerate
  
  localparam integer c0 = 0;
    generate 
        localparam integer d0 = 0;
        for (n0 = 0; n0 < 16; n0 = n0 + 1) 
        begin: outbit0
            assign data_11[n0 + d0*16 + c0*28*16] = data_11_array[c0][d0][n0];
        end
    endgenerate
    generate 
        localparam integer d1 = 1;
        for (n1 = 0; n1 < 16; n1 = n1 + 1) 
        begin: outbit1
            assign data_11[n1 + d1*16 + c0*28*16] = data_11_array[c0][d1][n1];
        end
    endgenerate
    generate 
        localparam integer d2 = 2;
        for (n2 = 0; n2 < 16; n2 = n2 + 1) 
        begin: outbit2
            assign data_11[n2 + d2*16 + c0*28*16] = data_11_array[c0][d2][n2];
        end
    endgenerate
    generate 
        localparam integer d3 = 3;
        for (n3 = 0; n3 < 16; n3 = n3 + 1) 
        begin: outbit3
            assign data_11[n3 + d3*16 + c0*28*16] = data_11_array[c0][d3][n3];
        end
    endgenerate
    generate 
        localparam integer d4 = 4;
        for (n4 = 0; n4 < 16; n4 = n4 + 1) 
        begin: outbit4
            assign data_11[n4 + d4*16 + c0*28*16] = data_11_array[c0][d4][n4];
        end
    endgenerate
    generate 
        localparam integer d5 = 5;
        for (n5 = 0; n5 < 16; n5 = n5 + 1) 
        begin: outbit5
            assign data_11[n5 + d5*16 + c0*28*16] = data_11_array[c0][d5][n5];
        end
    endgenerate
    generate 
        localparam integer d6 = 6;
        for (n6 = 0; n6 < 16; n6 = n6 + 1) 
        begin: outbit6
            assign data_11[n6 + d6*16 + c0*28*16] = data_11_array[c0][d6][n6];
        end
    endgenerate
    generate 
        localparam integer d7 = 7;
        for (n7 = 0; n7 < 16; n7 = n7 + 1) 
        begin: outbit7
            assign data_11[n7 + d7*16 + c0*28*16] = data_11_array[c0][d7][n7];
        end
    endgenerate
    generate 
        localparam integer d8 = 8;
        for (n8 = 0; n8 < 16; n8 = n8 + 1) 
        begin: outbit8
            assign data_11[n8 + d8*16 + c0*28*16] = data_11_array[c0][d8][n8];
        end
    endgenerate
    generate 
        localparam integer d9 = 9;
        for (n9 = 0; n9 < 16; n9 = n9 + 1) 
        begin: outbit9
            assign data_11[n9 + d9*16 + c0*28*16] = data_11_array[c0][d9][n9];
        end
    endgenerate
    generate 
        localparam integer d10 = 10;
        for (n10 = 0; n10 < 16; n10 = n10 + 1) 
        begin: outbit10
            assign data_11[n10 + d10*16 + c0*28*16] = data_11_array[c0][d10][n10];
        end
    endgenerate
    generate 
        localparam integer d11 = 11;
        for (n11 = 0; n11 < 16; n11 = n11 + 1) 
        begin: outbit11
            assign data_11[n11 + d11*16 + c0*28*16] = data_11_array[c0][d11][n11];
        end
    endgenerate
    generate 
        localparam integer d12 = 12;
        for (n12 = 0; n12 < 16; n12 = n12 + 1) 
        begin: outbit12
            assign data_11[n12 + d12*16 + c0*28*16] = data_11_array[c0][d12][n12];
        end
    endgenerate
    generate 
        localparam integer d13 = 13;
        for (n13 = 0; n13 < 16; n13 = n13 + 1) 
        begin: outbit13
            assign data_11[n13 + d13*16 + c0*28*16] = data_11_array[c0][d13][n13];
        end
    endgenerate
    generate 
        localparam integer d14 = 14;
        for (n14 = 0; n14 < 16; n14 = n14 + 1) 
        begin: outbit14
            assign data_11[n14 + d14*16 + c0*28*16] = data_11_array[c0][d14][n14];
        end
    endgenerate
    generate 
        localparam integer d15 = 15;
        for (n15 = 0; n15 < 16; n15 = n15 + 1) 
        begin: outbit15
            assign data_11[n15 + d15*16 + c0*28*16] = data_11_array[c0][d15][n15];
        end
    endgenerate
    generate 
        localparam integer d16 = 16;
        for (n16 = 0; n16 < 16; n16 = n16 + 1) 
        begin: outbit16
            assign data_11[n16 + d16*16 + c0*28*16] = data_11_array[c0][d16][n16];
        end
    endgenerate
    generate 
        localparam integer d17 = 17;
        for (n17 = 0; n17 < 16; n17 = n17 + 1) 
        begin: outbit17
            assign data_11[n17 + d17*16 + c0*28*16] = data_11_array[c0][d17][n17];
        end
    endgenerate
    generate 
        localparam integer d18 = 18;
        for (n18 = 0; n18 < 16; n18 = n18 + 1) 
        begin: outbit18
            assign data_11[n18 + d18*16 + c0*28*16] = data_11_array[c0][d18][n18];
        end
    endgenerate
    generate 
        localparam integer d19 = 19;
        for (n19 = 0; n19 < 16; n19 = n19 + 1) 
        begin: outbit19
            assign data_11[n19 + d19*16 + c0*28*16] = data_11_array[c0][d19][n19];
        end
    endgenerate
    generate 
        localparam integer d20 = 20;
        for (n20 = 0; n20 < 16; n20 = n20 + 1) 
        begin: outbit20
            assign data_11[n20 + d20*16 + c0*28*16] = data_11_array[c0][d20][n20];
        end
    endgenerate
    generate 
        localparam integer d21 = 21;
        for (n21 = 0; n21 < 16; n21 = n21 + 1) 
        begin: outbit21
            assign data_11[n21 + d21*16 + c0*28*16] = data_11_array[c0][d21][n21];
        end
    endgenerate
    generate 
        localparam integer d22 = 22;
        for (n22 = 0; n22 < 16; n22 = n22 + 1) 
        begin: outbit22
            assign data_11[n22 + d22*16 + c0*28*16] = data_11_array[c0][d22][n22];
        end
    endgenerate
    generate 
        localparam integer d23 = 23;
        for (n23 = 0; n23 < 16; n23 = n23 + 1) 
        begin: outbit23
            assign data_11[n23 + d23*16 + c0*28*16] = data_11_array[c0][d23][n23];
        end
    endgenerate
    generate 
        localparam integer d24 = 24;
        for (n24 = 0; n24 < 16; n24 = n24 + 1) 
        begin: outbit24
            assign data_11[n24 + d24*16 + c0*28*16] = data_11_array[c0][d24][n24];
        end
    endgenerate
    generate 
        localparam integer d25 = 25;
        for (n25 = 0; n25 < 16; n25 = n25 + 1) 
        begin: outbit25
            assign data_11[n25 + d25*16 + c0*28*16] = data_11_array[c0][d25][n25];
        end
    endgenerate
    generate 
        localparam integer d26 = 26;
        for (n26 = 0; n26 < 16; n26 = n26 + 1) 
        begin: outbit26
            assign data_11[n26 + d26*16 + c0*28*16] = data_11_array[c0][d26][n26];
        end
    endgenerate
    generate 
        localparam integer d27 = 27;
        for (n27 = 0; n27 < 16; n27 = n27 + 1) 
        begin: outbit27
            assign data_11[n27 + d27*16 + c0*28*16] = data_11_array[c0][d27][n27];
        end
    endgenerate
    localparam integer c1 = 1;
    generate 
        localparam integer d28 = 0;
        for (n28 = 0; n28 < 16; n28 = n28 + 1) 
        begin: outbit28
            assign data_11[n28 + d28*16 + c1*28*16] = data_11_array[c1][d28][n28];
        end
    endgenerate
    generate 
        localparam integer d29 = 1;
        for (n29 = 0; n29 < 16; n29 = n29 + 1) 
        begin: outbit29
            assign data_11[n29 + d29*16 + c1*28*16] = data_11_array[c1][d29][n29];
        end
    endgenerate
    generate 
        localparam integer d30 = 2;
        for (n30 = 0; n30 < 16; n30 = n30 + 1) 
        begin: outbit30
            assign data_11[n30 + d30*16 + c1*28*16] = data_11_array[c1][d30][n30];
        end
    endgenerate
    generate 
        localparam integer d31 = 3;
        for (n31 = 0; n31 < 16; n31 = n31 + 1) 
        begin: outbit31
            assign data_11[n31 + d31*16 + c1*28*16] = data_11_array[c1][d31][n31];
        end
    endgenerate
    generate 
        localparam integer d32 = 4;
        for (n32 = 0; n32 < 16; n32 = n32 + 1) 
        begin: outbit32
            assign data_11[n32 + d32*16 + c1*28*16] = data_11_array[c1][d32][n32];
        end
    endgenerate
    generate 
        localparam integer d33 = 5;
        for (n33 = 0; n33 < 16; n33 = n33 + 1) 
        begin: outbit33
            assign data_11[n33 + d33*16 + c1*28*16] = data_11_array[c1][d33][n33];
        end
    endgenerate
    generate 
        localparam integer d34 = 6;
        for (n34 = 0; n34 < 16; n34 = n34 + 1) 
        begin: outbit34
            assign data_11[n34 + d34*16 + c1*28*16] = data_11_array[c1][d34][n34];
        end
    endgenerate
    generate 
        localparam integer d35 = 7;
        for (n35 = 0; n35 < 16; n35 = n35 + 1) 
        begin: outbit35
            assign data_11[n35 + d35*16 + c1*28*16] = data_11_array[c1][d35][n35];
        end
    endgenerate
    generate 
        localparam integer d36 = 8;
        for (n36 = 0; n36 < 16; n36 = n36 + 1) 
        begin: outbit36
            assign data_11[n36 + d36*16 + c1*28*16] = data_11_array[c1][d36][n36];
        end
    endgenerate
    generate 
        localparam integer d37 = 9;
        for (n37 = 0; n37 < 16; n37 = n37 + 1) 
        begin: outbit37
            assign data_11[n37 + d37*16 + c1*28*16] = data_11_array[c1][d37][n37];
        end
    endgenerate
    generate 
        localparam integer d38 = 10;
        for (n38 = 0; n38 < 16; n38 = n38 + 1) 
        begin: outbit38
            assign data_11[n38 + d38*16 + c1*28*16] = data_11_array[c1][d38][n38];
        end
    endgenerate
    generate 
        localparam integer d39 = 11;
        for (n39 = 0; n39 < 16; n39 = n39 + 1) 
        begin: outbit39
            assign data_11[n39 + d39*16 + c1*28*16] = data_11_array[c1][d39][n39];
        end
    endgenerate
    generate 
        localparam integer d40 = 12;
        for (n40 = 0; n40 < 16; n40 = n40 + 1) 
        begin: outbit40
            assign data_11[n40 + d40*16 + c1*28*16] = data_11_array[c1][d40][n40];
        end
    endgenerate
    generate 
        localparam integer d41 = 13;
        for (n41 = 0; n41 < 16; n41 = n41 + 1) 
        begin: outbit41
            assign data_11[n41 + d41*16 + c1*28*16] = data_11_array[c1][d41][n41];
        end
    endgenerate
    generate 
        localparam integer d42 = 14;
        for (n42 = 0; n42 < 16; n42 = n42 + 1) 
        begin: outbit42
            assign data_11[n42 + d42*16 + c1*28*16] = data_11_array[c1][d42][n42];
        end
    endgenerate
    generate 
        localparam integer d43 = 15;
        for (n43 = 0; n43 < 16; n43 = n43 + 1) 
        begin: outbit43
            assign data_11[n43 + d43*16 + c1*28*16] = data_11_array[c1][d43][n43];
        end
    endgenerate
    generate 
        localparam integer d44 = 16;
        for (n44 = 0; n44 < 16; n44 = n44 + 1) 
        begin: outbit44
            assign data_11[n44 + d44*16 + c1*28*16] = data_11_array[c1][d44][n44];
        end
    endgenerate
    generate 
        localparam integer d45 = 17;
        for (n45 = 0; n45 < 16; n45 = n45 + 1) 
        begin: outbit45
            assign data_11[n45 + d45*16 + c1*28*16] = data_11_array[c1][d45][n45];
        end
    endgenerate
    generate 
        localparam integer d46 = 18;
        for (n46 = 0; n46 < 16; n46 = n46 + 1) 
        begin: outbit46
            assign data_11[n46 + d46*16 + c1*28*16] = data_11_array[c1][d46][n46];
        end
    endgenerate
    generate 
        localparam integer d47 = 19;
        for (n47 = 0; n47 < 16; n47 = n47 + 1) 
        begin: outbit47
            assign data_11[n47 + d47*16 + c1*28*16] = data_11_array[c1][d47][n47];
        end
    endgenerate
    generate 
        localparam integer d48 = 20;
        for (n48 = 0; n48 < 16; n48 = n48 + 1) 
        begin: outbit48
            assign data_11[n48 + d48*16 + c1*28*16] = data_11_array[c1][d48][n48];
        end
    endgenerate
    generate 
        localparam integer d49 = 21;
        for (n49 = 0; n49 < 16; n49 = n49 + 1) 
        begin: outbit49
            assign data_11[n49 + d49*16 + c1*28*16] = data_11_array[c1][d49][n49];
        end
    endgenerate
    generate 
        localparam integer d50 = 22;
        for (n50 = 0; n50 < 16; n50 = n50 + 1) 
        begin: outbit50
            assign data_11[n50 + d50*16 + c1*28*16] = data_11_array[c1][d50][n50];
        end
    endgenerate
    generate 
        localparam integer d51 = 23;
        for (n51 = 0; n51 < 16; n51 = n51 + 1) 
        begin: outbit51
            assign data_11[n51 + d51*16 + c1*28*16] = data_11_array[c1][d51][n51];
        end
    endgenerate
    generate 
        localparam integer d52 = 24;
        for (n52 = 0; n52 < 16; n52 = n52 + 1) 
        begin: outbit52
            assign data_11[n52 + d52*16 + c1*28*16] = data_11_array[c1][d52][n52];
        end
    endgenerate
    generate 
        localparam integer d53 = 25;
        for (n53 = 0; n53 < 16; n53 = n53 + 1) 
        begin: outbit53
            assign data_11[n53 + d53*16 + c1*28*16] = data_11_array[c1][d53][n53];
        end
    endgenerate
    generate 
        localparam integer d54 = 26;
        for (n54 = 0; n54 < 16; n54 = n54 + 1) 
        begin: outbit54
            assign data_11[n54 + d54*16 + c1*28*16] = data_11_array[c1][d54][n54];
        end
    endgenerate
    generate 
        localparam integer d55 = 27;
        for (n55 = 0; n55 < 16; n55 = n55 + 1) 
        begin: outbit55
            assign data_11[n55 + d55*16 + c1*28*16] = data_11_array[c1][d55][n55];
        end
    endgenerate
    localparam integer c2 = 2;
    generate 
        localparam integer d56 = 0;
        for (n56 = 0; n56 < 16; n56 = n56 + 1) 
        begin: outbit56
            assign data_11[n56 + d56*16 + c2*28*16] = data_11_array[c2][d56][n56];
        end
    endgenerate
    generate 
        localparam integer d57 = 1;
        for (n57 = 0; n57 < 16; n57 = n57 + 1) 
        begin: outbit57
            assign data_11[n57 + d57*16 + c2*28*16] = data_11_array[c2][d57][n57];
        end
    endgenerate
    generate 
        localparam integer d58 = 2;
        for (n58 = 0; n58 < 16; n58 = n58 + 1) 
        begin: outbit58
            assign data_11[n58 + d58*16 + c2*28*16] = data_11_array[c2][d58][n58];
        end
    endgenerate
    generate 
        localparam integer d59 = 3;
        for (n59 = 0; n59 < 16; n59 = n59 + 1) 
        begin: outbit59
            assign data_11[n59 + d59*16 + c2*28*16] = data_11_array[c2][d59][n59];
        end
    endgenerate
    generate 
        localparam integer d60 = 4;
        for (n60 = 0; n60 < 16; n60 = n60 + 1) 
        begin: outbit60
            assign data_11[n60 + d60*16 + c2*28*16] = data_11_array[c2][d60][n60];
        end
    endgenerate
    generate 
        localparam integer d61 = 5;
        for (n61 = 0; n61 < 16; n61 = n61 + 1) 
        begin: outbit61
            assign data_11[n61 + d61*16 + c2*28*16] = data_11_array[c2][d61][n61];
        end
    endgenerate
    generate 
        localparam integer d62 = 6;
        for (n62 = 0; n62 < 16; n62 = n62 + 1) 
        begin: outbit62
            assign data_11[n62 + d62*16 + c2*28*16] = data_11_array[c2][d62][n62];
        end
    endgenerate
    generate 
        localparam integer d63 = 7;
        for (n63 = 0; n63 < 16; n63 = n63 + 1) 
        begin: outbit63
            assign data_11[n63 + d63*16 + c2*28*16] = data_11_array[c2][d63][n63];
        end
    endgenerate
    generate 
        localparam integer d64 = 8;
        for (n64 = 0; n64 < 16; n64 = n64 + 1) 
        begin: outbit64
            assign data_11[n64 + d64*16 + c2*28*16] = data_11_array[c2][d64][n64];
        end
    endgenerate
    generate 
        localparam integer d65 = 9;
        for (n65 = 0; n65 < 16; n65 = n65 + 1) 
        begin: outbit65
            assign data_11[n65 + d65*16 + c2*28*16] = data_11_array[c2][d65][n65];
        end
    endgenerate
    generate 
        localparam integer d66 = 10;
        for (n66 = 0; n66 < 16; n66 = n66 + 1) 
        begin: outbit66
            assign data_11[n66 + d66*16 + c2*28*16] = data_11_array[c2][d66][n66];
        end
    endgenerate
    generate 
        localparam integer d67 = 11;
        for (n67 = 0; n67 < 16; n67 = n67 + 1) 
        begin: outbit67
            assign data_11[n67 + d67*16 + c2*28*16] = data_11_array[c2][d67][n67];
        end
    endgenerate
    generate 
        localparam integer d68 = 12;
        for (n68 = 0; n68 < 16; n68 = n68 + 1) 
        begin: outbit68
            assign data_11[n68 + d68*16 + c2*28*16] = data_11_array[c2][d68][n68];
        end
    endgenerate
    generate 
        localparam integer d69 = 13;
        for (n69 = 0; n69 < 16; n69 = n69 + 1) 
        begin: outbit69
            assign data_11[n69 + d69*16 + c2*28*16] = data_11_array[c2][d69][n69];
        end
    endgenerate
    generate 
        localparam integer d70 = 14;
        for (n70 = 0; n70 < 16; n70 = n70 + 1) 
        begin: outbit70
            assign data_11[n70 + d70*16 + c2*28*16] = data_11_array[c2][d70][n70];
        end
    endgenerate
    generate 
        localparam integer d71 = 15;
        for (n71 = 0; n71 < 16; n71 = n71 + 1) 
        begin: outbit71
            assign data_11[n71 + d71*16 + c2*28*16] = data_11_array[c2][d71][n71];
        end
    endgenerate
    generate 
        localparam integer d72 = 16;
        for (n72 = 0; n72 < 16; n72 = n72 + 1) 
        begin: outbit72
            assign data_11[n72 + d72*16 + c2*28*16] = data_11_array[c2][d72][n72];
        end
    endgenerate
    generate 
        localparam integer d73 = 17;
        for (n73 = 0; n73 < 16; n73 = n73 + 1) 
        begin: outbit73
            assign data_11[n73 + d73*16 + c2*28*16] = data_11_array[c2][d73][n73];
        end
    endgenerate
    generate 
        localparam integer d74 = 18;
        for (n74 = 0; n74 < 16; n74 = n74 + 1) 
        begin: outbit74
            assign data_11[n74 + d74*16 + c2*28*16] = data_11_array[c2][d74][n74];
        end
    endgenerate
    generate 
        localparam integer d75 = 19;
        for (n75 = 0; n75 < 16; n75 = n75 + 1) 
        begin: outbit75
            assign data_11[n75 + d75*16 + c2*28*16] = data_11_array[c2][d75][n75];
        end
    endgenerate
    generate 
        localparam integer d76 = 20;
        for (n76 = 0; n76 < 16; n76 = n76 + 1) 
        begin: outbit76
            assign data_11[n76 + d76*16 + c2*28*16] = data_11_array[c2][d76][n76];
        end
    endgenerate
    generate 
        localparam integer d77 = 21;
        for (n77 = 0; n77 < 16; n77 = n77 + 1) 
        begin: outbit77
            assign data_11[n77 + d77*16 + c2*28*16] = data_11_array[c2][d77][n77];
        end
    endgenerate
    generate 
        localparam integer d78 = 22;
        for (n78 = 0; n78 < 16; n78 = n78 + 1) 
        begin: outbit78
            assign data_11[n78 + d78*16 + c2*28*16] = data_11_array[c2][d78][n78];
        end
    endgenerate
    generate 
        localparam integer d79 = 23;
        for (n79 = 0; n79 < 16; n79 = n79 + 1) 
        begin: outbit79
            assign data_11[n79 + d79*16 + c2*28*16] = data_11_array[c2][d79][n79];
        end
    endgenerate
    generate 
        localparam integer d80 = 24;
        for (n80 = 0; n80 < 16; n80 = n80 + 1) 
        begin: outbit80
            assign data_11[n80 + d80*16 + c2*28*16] = data_11_array[c2][d80][n80];
        end
    endgenerate
    generate 
        localparam integer d81 = 25;
        for (n81 = 0; n81 < 16; n81 = n81 + 1) 
        begin: outbit81
            assign data_11[n81 + d81*16 + c2*28*16] = data_11_array[c2][d81][n81];
        end
    endgenerate
    generate 
        localparam integer d82 = 26;
        for (n82 = 0; n82 < 16; n82 = n82 + 1) 
        begin: outbit82
            assign data_11[n82 + d82*16 + c2*28*16] = data_11_array[c2][d82][n82];
        end
    endgenerate
    generate 
        localparam integer d83 = 27;
        for (n83 = 0; n83 < 16; n83 = n83 + 1) 
        begin: outbit83
            assign data_11[n83 + d83*16 + c2*28*16] = data_11_array[c2][d83][n83];
        end
    endgenerate
    localparam integer c3 = 3;
    generate 
        localparam integer d84 = 0;
        for (n84 = 0; n84 < 16; n84 = n84 + 1) 
        begin: outbit84
            assign data_11[n84 + d84*16 + c3*28*16] = data_11_array[c3][d84][n84];
        end
    endgenerate
    generate 
        localparam integer d85 = 1;
        for (n85 = 0; n85 < 16; n85 = n85 + 1) 
        begin: outbit85
            assign data_11[n85 + d85*16 + c3*28*16] = data_11_array[c3][d85][n85];
        end
    endgenerate
    generate 
        localparam integer d86 = 2;
        for (n86 = 0; n86 < 16; n86 = n86 + 1) 
        begin: outbit86
            assign data_11[n86 + d86*16 + c3*28*16] = data_11_array[c3][d86][n86];
        end
    endgenerate
    generate 
        localparam integer d87 = 3;
        for (n87 = 0; n87 < 16; n87 = n87 + 1) 
        begin: outbit87
            assign data_11[n87 + d87*16 + c3*28*16] = data_11_array[c3][d87][n87];
        end
    endgenerate
    generate 
        localparam integer d88 = 4;
        for (n88 = 0; n88 < 16; n88 = n88 + 1) 
        begin: outbit88
            assign data_11[n88 + d88*16 + c3*28*16] = data_11_array[c3][d88][n88];
        end
    endgenerate
    generate 
        localparam integer d89 = 5;
        for (n89 = 0; n89 < 16; n89 = n89 + 1) 
        begin: outbit89
            assign data_11[n89 + d89*16 + c3*28*16] = data_11_array[c3][d89][n89];
        end
    endgenerate
    generate 
        localparam integer d90 = 6;
        for (n90 = 0; n90 < 16; n90 = n90 + 1) 
        begin: outbit90
            assign data_11[n90 + d90*16 + c3*28*16] = data_11_array[c3][d90][n90];
        end
    endgenerate
    generate 
        localparam integer d91 = 7;
        for (n91 = 0; n91 < 16; n91 = n91 + 1) 
        begin: outbit91
            assign data_11[n91 + d91*16 + c3*28*16] = data_11_array[c3][d91][n91];
        end
    endgenerate
    generate 
        localparam integer d92 = 8;
        for (n92 = 0; n92 < 16; n92 = n92 + 1) 
        begin: outbit92
            assign data_11[n92 + d92*16 + c3*28*16] = data_11_array[c3][d92][n92];
        end
    endgenerate
    generate 
        localparam integer d93 = 9;
        for (n93 = 0; n93 < 16; n93 = n93 + 1) 
        begin: outbit93
            assign data_11[n93 + d93*16 + c3*28*16] = data_11_array[c3][d93][n93];
        end
    endgenerate
    generate 
        localparam integer d94 = 10;
        for (n94 = 0; n94 < 16; n94 = n94 + 1) 
        begin: outbit94
            assign data_11[n94 + d94*16 + c3*28*16] = data_11_array[c3][d94][n94];
        end
    endgenerate
    generate 
        localparam integer d95 = 11;
        for (n95 = 0; n95 < 16; n95 = n95 + 1) 
        begin: outbit95
            assign data_11[n95 + d95*16 + c3*28*16] = data_11_array[c3][d95][n95];
        end
    endgenerate
    generate 
        localparam integer d96 = 12;
        for (n96 = 0; n96 < 16; n96 = n96 + 1) 
        begin: outbit96
            assign data_11[n96 + d96*16 + c3*28*16] = data_11_array[c3][d96][n96];
        end
    endgenerate
    generate 
        localparam integer d97 = 13;
        for (n97 = 0; n97 < 16; n97 = n97 + 1) 
        begin: outbit97
            assign data_11[n97 + d97*16 + c3*28*16] = data_11_array[c3][d97][n97];
        end
    endgenerate
    generate 
        localparam integer d98 = 14;
        for (n98 = 0; n98 < 16; n98 = n98 + 1) 
        begin: outbit98
            assign data_11[n98 + d98*16 + c3*28*16] = data_11_array[c3][d98][n98];
        end
    endgenerate
    generate 
        localparam integer d99 = 15;
        for (n99 = 0; n99 < 16; n99 = n99 + 1) 
        begin: outbit99
            assign data_11[n99 + d99*16 + c3*28*16] = data_11_array[c3][d99][n99];
        end
    endgenerate
    generate 
        localparam integer d100 = 16;
        for (n100 = 0; n100 < 16; n100 = n100 + 1) 
        begin: outbit100
            assign data_11[n100 + d100*16 + c3*28*16] = data_11_array[c3][d100][n100];
        end
    endgenerate
    generate 
        localparam integer d101 = 17;
        for (n101 = 0; n101 < 16; n101 = n101 + 1) 
        begin: outbit101
            assign data_11[n101 + d101*16 + c3*28*16] = data_11_array[c3][d101][n101];
        end
    endgenerate
    generate 
        localparam integer d102 = 18;
        for (n102 = 0; n102 < 16; n102 = n102 + 1) 
        begin: outbit102
            assign data_11[n102 + d102*16 + c3*28*16] = data_11_array[c3][d102][n102];
        end
    endgenerate
    generate 
        localparam integer d103 = 19;
        for (n103 = 0; n103 < 16; n103 = n103 + 1) 
        begin: outbit103
            assign data_11[n103 + d103*16 + c3*28*16] = data_11_array[c3][d103][n103];
        end
    endgenerate
    generate 
        localparam integer d104 = 20;
        for (n104 = 0; n104 < 16; n104 = n104 + 1) 
        begin: outbit104
            assign data_11[n104 + d104*16 + c3*28*16] = data_11_array[c3][d104][n104];
        end
    endgenerate
    generate 
        localparam integer d105 = 21;
        for (n105 = 0; n105 < 16; n105 = n105 + 1) 
        begin: outbit105
            assign data_11[n105 + d105*16 + c3*28*16] = data_11_array[c3][d105][n105];
        end
    endgenerate
    generate 
        localparam integer d106 = 22;
        for (n106 = 0; n106 < 16; n106 = n106 + 1) 
        begin: outbit106
            assign data_11[n106 + d106*16 + c3*28*16] = data_11_array[c3][d106][n106];
        end
    endgenerate
    generate 
        localparam integer d107 = 23;
        for (n107 = 0; n107 < 16; n107 = n107 + 1) 
        begin: outbit107
            assign data_11[n107 + d107*16 + c3*28*16] = data_11_array[c3][d107][n107];
        end
    endgenerate
    generate 
        localparam integer d108 = 24;
        for (n108 = 0; n108 < 16; n108 = n108 + 1) 
        begin: outbit108
            assign data_11[n108 + d108*16 + c3*28*16] = data_11_array[c3][d108][n108];
        end
    endgenerate
    generate 
        localparam integer d109 = 25;
        for (n109 = 0; n109 < 16; n109 = n109 + 1) 
        begin: outbit109
            assign data_11[n109 + d109*16 + c3*28*16] = data_11_array[c3][d109][n109];
        end
    endgenerate
    generate 
        localparam integer d110 = 26;
        for (n110 = 0; n110 < 16; n110 = n110 + 1) 
        begin: outbit110
            assign data_11[n110 + d110*16 + c3*28*16] = data_11_array[c3][d110][n110];
        end
    endgenerate
    generate 
        localparam integer d111 = 27;
        for (n111 = 0; n111 < 16; n111 = n111 + 1) 
        begin: outbit111
            assign data_11[n111 + d111*16 + c3*28*16] = data_11_array[c3][d111][n111];
        end
    endgenerate
    localparam integer c4 = 4;
    generate 
        localparam integer d112 = 0;
        for (n112 = 0; n112 < 16; n112 = n112 + 1) 
        begin: outbit112
            assign data_11[n112 + d112*16 + c4*28*16] = data_11_array[c4][d112][n112];
        end
    endgenerate
    generate 
        localparam integer d113 = 1;
        for (n113 = 0; n113 < 16; n113 = n113 + 1) 
        begin: outbit113
            assign data_11[n113 + d113*16 + c4*28*16] = data_11_array[c4][d113][n113];
        end
    endgenerate
    generate 
        localparam integer d114 = 2;
        for (n114 = 0; n114 < 16; n114 = n114 + 1) 
        begin: outbit114
            assign data_11[n114 + d114*16 + c4*28*16] = data_11_array[c4][d114][n114];
        end
    endgenerate
    generate 
        localparam integer d115 = 3;
        for (n115 = 0; n115 < 16; n115 = n115 + 1) 
        begin: outbit115
            assign data_11[n115 + d115*16 + c4*28*16] = data_11_array[c4][d115][n115];
        end
    endgenerate
    generate 
        localparam integer d116 = 4;
        for (n116 = 0; n116 < 16; n116 = n116 + 1) 
        begin: outbit116
            assign data_11[n116 + d116*16 + c4*28*16] = data_11_array[c4][d116][n116];
        end
    endgenerate
    generate 
        localparam integer d117 = 5;
        for (n117 = 0; n117 < 16; n117 = n117 + 1) 
        begin: outbit117
            assign data_11[n117 + d117*16 + c4*28*16] = data_11_array[c4][d117][n117];
        end
    endgenerate
    generate 
        localparam integer d118 = 6;
        for (n118 = 0; n118 < 16; n118 = n118 + 1) 
        begin: outbit118
            assign data_11[n118 + d118*16 + c4*28*16] = data_11_array[c4][d118][n118];
        end
    endgenerate
    generate 
        localparam integer d119 = 7;
        for (n119 = 0; n119 < 16; n119 = n119 + 1) 
        begin: outbit119
            assign data_11[n119 + d119*16 + c4*28*16] = data_11_array[c4][d119][n119];
        end
    endgenerate
    generate 
        localparam integer d120 = 8;
        for (n120 = 0; n120 < 16; n120 = n120 + 1) 
        begin: outbit120
            assign data_11[n120 + d120*16 + c4*28*16] = data_11_array[c4][d120][n120];
        end
    endgenerate
    generate 
        localparam integer d121 = 9;
        for (n121 = 0; n121 < 16; n121 = n121 + 1) 
        begin: outbit121
            assign data_11[n121 + d121*16 + c4*28*16] = data_11_array[c4][d121][n121];
        end
    endgenerate
    generate 
        localparam integer d122 = 10;
        for (n122 = 0; n122 < 16; n122 = n122 + 1) 
        begin: outbit122
            assign data_11[n122 + d122*16 + c4*28*16] = data_11_array[c4][d122][n122];
        end
    endgenerate
    generate 
        localparam integer d123 = 11;
        for (n123 = 0; n123 < 16; n123 = n123 + 1) 
        begin: outbit123
            assign data_11[n123 + d123*16 + c4*28*16] = data_11_array[c4][d123][n123];
        end
    endgenerate
    generate 
        localparam integer d124 = 12;
        for (n124 = 0; n124 < 16; n124 = n124 + 1) 
        begin: outbit124
            assign data_11[n124 + d124*16 + c4*28*16] = data_11_array[c4][d124][n124];
        end
    endgenerate
    generate 
        localparam integer d125 = 13;
        for (n125 = 0; n125 < 16; n125 = n125 + 1) 
        begin: outbit125
            assign data_11[n125 + d125*16 + c4*28*16] = data_11_array[c4][d125][n125];
        end
    endgenerate
    generate 
        localparam integer d126 = 14;
        for (n126 = 0; n126 < 16; n126 = n126 + 1) 
        begin: outbit126
            assign data_11[n126 + d126*16 + c4*28*16] = data_11_array[c4][d126][n126];
        end
    endgenerate
    generate 
        localparam integer d127 = 15;
        for (n127 = 0; n127 < 16; n127 = n127 + 1) 
        begin: outbit127
            assign data_11[n127 + d127*16 + c4*28*16] = data_11_array[c4][d127][n127];
        end
    endgenerate
    generate 
        localparam integer d128 = 16;
        for (n128 = 0; n128 < 16; n128 = n128 + 1) 
        begin: outbit128
            assign data_11[n128 + d128*16 + c4*28*16] = data_11_array[c4][d128][n128];
        end
    endgenerate
    generate 
        localparam integer d129 = 17;
        for (n129 = 0; n129 < 16; n129 = n129 + 1) 
        begin: outbit129
            assign data_11[n129 + d129*16 + c4*28*16] = data_11_array[c4][d129][n129];
        end
    endgenerate
    generate 
        localparam integer d130 = 18;
        for (n130 = 0; n130 < 16; n130 = n130 + 1) 
        begin: outbit130
            assign data_11[n130 + d130*16 + c4*28*16] = data_11_array[c4][d130][n130];
        end
    endgenerate
    generate 
        localparam integer d131 = 19;
        for (n131 = 0; n131 < 16; n131 = n131 + 1) 
        begin: outbit131
            assign data_11[n131 + d131*16 + c4*28*16] = data_11_array[c4][d131][n131];
        end
    endgenerate
    generate 
        localparam integer d132 = 20;
        for (n132 = 0; n132 < 16; n132 = n132 + 1) 
        begin: outbit132
            assign data_11[n132 + d132*16 + c4*28*16] = data_11_array[c4][d132][n132];
        end
    endgenerate
    generate 
        localparam integer d133 = 21;
        for (n133 = 0; n133 < 16; n133 = n133 + 1) 
        begin: outbit133
            assign data_11[n133 + d133*16 + c4*28*16] = data_11_array[c4][d133][n133];
        end
    endgenerate
    generate 
        localparam integer d134 = 22;
        for (n134 = 0; n134 < 16; n134 = n134 + 1) 
        begin: outbit134
            assign data_11[n134 + d134*16 + c4*28*16] = data_11_array[c4][d134][n134];
        end
    endgenerate
    generate 
        localparam integer d135 = 23;
        for (n135 = 0; n135 < 16; n135 = n135 + 1) 
        begin: outbit135
            assign data_11[n135 + d135*16 + c4*28*16] = data_11_array[c4][d135][n135];
        end
    endgenerate
    generate 
        localparam integer d136 = 24;
        for (n136 = 0; n136 < 16; n136 = n136 + 1) 
        begin: outbit136
            assign data_11[n136 + d136*16 + c4*28*16] = data_11_array[c4][d136][n136];
        end
    endgenerate
    generate 
        localparam integer d137 = 25;
        for (n137 = 0; n137 < 16; n137 = n137 + 1) 
        begin: outbit137
            assign data_11[n137 + d137*16 + c4*28*16] = data_11_array[c4][d137][n137];
        end
    endgenerate
    generate 
        localparam integer d138 = 26;
        for (n138 = 0; n138 < 16; n138 = n138 + 1) 
        begin: outbit138
            assign data_11[n138 + d138*16 + c4*28*16] = data_11_array[c4][d138][n138];
        end
    endgenerate
    generate 
        localparam integer d139 = 27;
        for (n139 = 0; n139 < 16; n139 = n139 + 1) 
        begin: outbit139
            assign data_11[n139 + d139*16 + c4*28*16] = data_11_array[c4][d139][n139];
        end
    endgenerate
    localparam integer c5 = 5;
    generate 
        localparam integer d140 = 0;
        for (n140 = 0; n140 < 16; n140 = n140 + 1) 
        begin: outbit140
            assign data_11[n140 + d140*16 + c5*28*16] = data_11_array[c5][d140][n140];
        end
    endgenerate
    generate 
        localparam integer d141 = 1;
        for (n141 = 0; n141 < 16; n141 = n141 + 1) 
        begin: outbit141
            assign data_11[n141 + d141*16 + c5*28*16] = data_11_array[c5][d141][n141];
        end
    endgenerate
    generate 
        localparam integer d142 = 2;
        for (n142 = 0; n142 < 16; n142 = n142 + 1) 
        begin: outbit142
            assign data_11[n142 + d142*16 + c5*28*16] = data_11_array[c5][d142][n142];
        end
    endgenerate
    generate 
        localparam integer d143 = 3;
        for (n143 = 0; n143 < 16; n143 = n143 + 1) 
        begin: outbit143
            assign data_11[n143 + d143*16 + c5*28*16] = data_11_array[c5][d143][n143];
        end
    endgenerate
    generate 
        localparam integer d144 = 4;
        for (n144 = 0; n144 < 16; n144 = n144 + 1) 
        begin: outbit144
            assign data_11[n144 + d144*16 + c5*28*16] = data_11_array[c5][d144][n144];
        end
    endgenerate
    generate 
        localparam integer d145 = 5;
        for (n145 = 0; n145 < 16; n145 = n145 + 1) 
        begin: outbit145
            assign data_11[n145 + d145*16 + c5*28*16] = data_11_array[c5][d145][n145];
        end
    endgenerate
    generate 
        localparam integer d146 = 6;
        for (n146 = 0; n146 < 16; n146 = n146 + 1) 
        begin: outbit146
            assign data_11[n146 + d146*16 + c5*28*16] = data_11_array[c5][d146][n146];
        end
    endgenerate
    generate 
        localparam integer d147 = 7;
        for (n147 = 0; n147 < 16; n147 = n147 + 1) 
        begin: outbit147
            assign data_11[n147 + d147*16 + c5*28*16] = data_11_array[c5][d147][n147];
        end
    endgenerate
    generate 
        localparam integer d148 = 8;
        for (n148 = 0; n148 < 16; n148 = n148 + 1) 
        begin: outbit148
            assign data_11[n148 + d148*16 + c5*28*16] = data_11_array[c5][d148][n148];
        end
    endgenerate
    generate 
        localparam integer d149 = 9;
        for (n149 = 0; n149 < 16; n149 = n149 + 1) 
        begin: outbit149
            assign data_11[n149 + d149*16 + c5*28*16] = data_11_array[c5][d149][n149];
        end
    endgenerate
    generate 
        localparam integer d150 = 10;
        for (n150 = 0; n150 < 16; n150 = n150 + 1) 
        begin: outbit150
            assign data_11[n150 + d150*16 + c5*28*16] = data_11_array[c5][d150][n150];
        end
    endgenerate
    generate 
        localparam integer d151 = 11;
        for (n151 = 0; n151 < 16; n151 = n151 + 1) 
        begin: outbit151
            assign data_11[n151 + d151*16 + c5*28*16] = data_11_array[c5][d151][n151];
        end
    endgenerate
    generate 
        localparam integer d152 = 12;
        for (n152 = 0; n152 < 16; n152 = n152 + 1) 
        begin: outbit152
            assign data_11[n152 + d152*16 + c5*28*16] = data_11_array[c5][d152][n152];
        end
    endgenerate
    generate 
        localparam integer d153 = 13;
        for (n153 = 0; n153 < 16; n153 = n153 + 1) 
        begin: outbit153
            assign data_11[n153 + d153*16 + c5*28*16] = data_11_array[c5][d153][n153];
        end
    endgenerate
    generate 
        localparam integer d154 = 14;
        for (n154 = 0; n154 < 16; n154 = n154 + 1) 
        begin: outbit154
            assign data_11[n154 + d154*16 + c5*28*16] = data_11_array[c5][d154][n154];
        end
    endgenerate
    generate 
        localparam integer d155 = 15;
        for (n155 = 0; n155 < 16; n155 = n155 + 1) 
        begin: outbit155
            assign data_11[n155 + d155*16 + c5*28*16] = data_11_array[c5][d155][n155];
        end
    endgenerate
    generate 
        localparam integer d156 = 16;
        for (n156 = 0; n156 < 16; n156 = n156 + 1) 
        begin: outbit156
            assign data_11[n156 + d156*16 + c5*28*16] = data_11_array[c5][d156][n156];
        end
    endgenerate
    generate 
        localparam integer d157 = 17;
        for (n157 = 0; n157 < 16; n157 = n157 + 1) 
        begin: outbit157
            assign data_11[n157 + d157*16 + c5*28*16] = data_11_array[c5][d157][n157];
        end
    endgenerate
    generate 
        localparam integer d158 = 18;
        for (n158 = 0; n158 < 16; n158 = n158 + 1) 
        begin: outbit158
            assign data_11[n158 + d158*16 + c5*28*16] = data_11_array[c5][d158][n158];
        end
    endgenerate
    generate 
        localparam integer d159 = 19;
        for (n159 = 0; n159 < 16; n159 = n159 + 1) 
        begin: outbit159
            assign data_11[n159 + d159*16 + c5*28*16] = data_11_array[c5][d159][n159];
        end
    endgenerate
    generate 
        localparam integer d160 = 20;
        for (n160 = 0; n160 < 16; n160 = n160 + 1) 
        begin: outbit160
            assign data_11[n160 + d160*16 + c5*28*16] = data_11_array[c5][d160][n160];
        end
    endgenerate
    generate 
        localparam integer d161 = 21;
        for (n161 = 0; n161 < 16; n161 = n161 + 1) 
        begin: outbit161
            assign data_11[n161 + d161*16 + c5*28*16] = data_11_array[c5][d161][n161];
        end
    endgenerate
    generate 
        localparam integer d162 = 22;
        for (n162 = 0; n162 < 16; n162 = n162 + 1) 
        begin: outbit162
            assign data_11[n162 + d162*16 + c5*28*16] = data_11_array[c5][d162][n162];
        end
    endgenerate
    generate 
        localparam integer d163 = 23;
        for (n163 = 0; n163 < 16; n163 = n163 + 1) 
        begin: outbit163
            assign data_11[n163 + d163*16 + c5*28*16] = data_11_array[c5][d163][n163];
        end
    endgenerate
    generate 
        localparam integer d164 = 24;
        for (n164 = 0; n164 < 16; n164 = n164 + 1) 
        begin: outbit164
            assign data_11[n164 + d164*16 + c5*28*16] = data_11_array[c5][d164][n164];
        end
    endgenerate
    generate 
        localparam integer d165 = 25;
        for (n165 = 0; n165 < 16; n165 = n165 + 1) 
        begin: outbit165
            assign data_11[n165 + d165*16 + c5*28*16] = data_11_array[c5][d165][n165];
        end
    endgenerate
    generate 
        localparam integer d166 = 26;
        for (n166 = 0; n166 < 16; n166 = n166 + 1) 
        begin: outbit166
            assign data_11[n166 + d166*16 + c5*28*16] = data_11_array[c5][d166][n166];
        end
    endgenerate
    generate 
        localparam integer d167 = 27;
        for (n167 = 0; n167 < 16; n167 = n167 + 1) 
        begin: outbit167
            assign data_11[n167 + d167*16 + c5*28*16] = data_11_array[c5][d167][n167];
        end
    endgenerate
    localparam integer c6 = 6;
    generate 
        localparam integer d168 = 0;
        for (n168 = 0; n168 < 16; n168 = n168 + 1) 
        begin: outbit168
            assign data_11[n168 + d168*16 + c6*28*16] = data_11_array[c6][d168][n168];
        end
    endgenerate
    generate 
        localparam integer d169 = 1;
        for (n169 = 0; n169 < 16; n169 = n169 + 1) 
        begin: outbit169
            assign data_11[n169 + d169*16 + c6*28*16] = data_11_array[c6][d169][n169];
        end
    endgenerate
    generate 
        localparam integer d170 = 2;
        for (n170 = 0; n170 < 16; n170 = n170 + 1) 
        begin: outbit170
            assign data_11[n170 + d170*16 + c6*28*16] = data_11_array[c6][d170][n170];
        end
    endgenerate
    generate 
        localparam integer d171 = 3;
        for (n171 = 0; n171 < 16; n171 = n171 + 1) 
        begin: outbit171
            assign data_11[n171 + d171*16 + c6*28*16] = data_11_array[c6][d171][n171];
        end
    endgenerate
    generate 
        localparam integer d172 = 4;
        for (n172 = 0; n172 < 16; n172 = n172 + 1) 
        begin: outbit172
            assign data_11[n172 + d172*16 + c6*28*16] = data_11_array[c6][d172][n172];
        end
    endgenerate
    generate 
        localparam integer d173 = 5;
        for (n173 = 0; n173 < 16; n173 = n173 + 1) 
        begin: outbit173
            assign data_11[n173 + d173*16 + c6*28*16] = data_11_array[c6][d173][n173];
        end
    endgenerate
    generate 
        localparam integer d174 = 6;
        for (n174 = 0; n174 < 16; n174 = n174 + 1) 
        begin: outbit174
            assign data_11[n174 + d174*16 + c6*28*16] = data_11_array[c6][d174][n174];
        end
    endgenerate
    generate 
        localparam integer d175 = 7;
        for (n175 = 0; n175 < 16; n175 = n175 + 1) 
        begin: outbit175
            assign data_11[n175 + d175*16 + c6*28*16] = data_11_array[c6][d175][n175];
        end
    endgenerate
    generate 
        localparam integer d176 = 8;
        for (n176 = 0; n176 < 16; n176 = n176 + 1) 
        begin: outbit176
            assign data_11[n176 + d176*16 + c6*28*16] = data_11_array[c6][d176][n176];
        end
    endgenerate
    generate 
        localparam integer d177 = 9;
        for (n177 = 0; n177 < 16; n177 = n177 + 1) 
        begin: outbit177
            assign data_11[n177 + d177*16 + c6*28*16] = data_11_array[c6][d177][n177];
        end
    endgenerate
    generate 
        localparam integer d178 = 10;
        for (n178 = 0; n178 < 16; n178 = n178 + 1) 
        begin: outbit178
            assign data_11[n178 + d178*16 + c6*28*16] = data_11_array[c6][d178][n178];
        end
    endgenerate
    generate 
        localparam integer d179 = 11;
        for (n179 = 0; n179 < 16; n179 = n179 + 1) 
        begin: outbit179
            assign data_11[n179 + d179*16 + c6*28*16] = data_11_array[c6][d179][n179];
        end
    endgenerate
    generate 
        localparam integer d180 = 12;
        for (n180 = 0; n180 < 16; n180 = n180 + 1) 
        begin: outbit180
            assign data_11[n180 + d180*16 + c6*28*16] = data_11_array[c6][d180][n180];
        end
    endgenerate
    generate 
        localparam integer d181 = 13;
        for (n181 = 0; n181 < 16; n181 = n181 + 1) 
        begin: outbit181
            assign data_11[n181 + d181*16 + c6*28*16] = data_11_array[c6][d181][n181];
        end
    endgenerate
    generate 
        localparam integer d182 = 14;
        for (n182 = 0; n182 < 16; n182 = n182 + 1) 
        begin: outbit182
            assign data_11[n182 + d182*16 + c6*28*16] = data_11_array[c6][d182][n182];
        end
    endgenerate
    generate 
        localparam integer d183 = 15;
        for (n183 = 0; n183 < 16; n183 = n183 + 1) 
        begin: outbit183
            assign data_11[n183 + d183*16 + c6*28*16] = data_11_array[c6][d183][n183];
        end
    endgenerate
    generate 
        localparam integer d184 = 16;
        for (n184 = 0; n184 < 16; n184 = n184 + 1) 
        begin: outbit184
            assign data_11[n184 + d184*16 + c6*28*16] = data_11_array[c6][d184][n184];
        end
    endgenerate
    generate 
        localparam integer d185 = 17;
        for (n185 = 0; n185 < 16; n185 = n185 + 1) 
        begin: outbit185
            assign data_11[n185 + d185*16 + c6*28*16] = data_11_array[c6][d185][n185];
        end
    endgenerate
    generate 
        localparam integer d186 = 18;
        for (n186 = 0; n186 < 16; n186 = n186 + 1) 
        begin: outbit186
            assign data_11[n186 + d186*16 + c6*28*16] = data_11_array[c6][d186][n186];
        end
    endgenerate
    generate 
        localparam integer d187 = 19;
        for (n187 = 0; n187 < 16; n187 = n187 + 1) 
        begin: outbit187
            assign data_11[n187 + d187*16 + c6*28*16] = data_11_array[c6][d187][n187];
        end
    endgenerate
    generate 
        localparam integer d188 = 20;
        for (n188 = 0; n188 < 16; n188 = n188 + 1) 
        begin: outbit188
            assign data_11[n188 + d188*16 + c6*28*16] = data_11_array[c6][d188][n188];
        end
    endgenerate
    generate 
        localparam integer d189 = 21;
        for (n189 = 0; n189 < 16; n189 = n189 + 1) 
        begin: outbit189
            assign data_11[n189 + d189*16 + c6*28*16] = data_11_array[c6][d189][n189];
        end
    endgenerate
    generate 
        localparam integer d190 = 22;
        for (n190 = 0; n190 < 16; n190 = n190 + 1) 
        begin: outbit190
            assign data_11[n190 + d190*16 + c6*28*16] = data_11_array[c6][d190][n190];
        end
    endgenerate
    generate 
        localparam integer d191 = 23;
        for (n191 = 0; n191 < 16; n191 = n191 + 1) 
        begin: outbit191
            assign data_11[n191 + d191*16 + c6*28*16] = data_11_array[c6][d191][n191];
        end
    endgenerate
    generate 
        localparam integer d192 = 24;
        for (n192 = 0; n192 < 16; n192 = n192 + 1) 
        begin: outbit192
            assign data_11[n192 + d192*16 + c6*28*16] = data_11_array[c6][d192][n192];
        end
    endgenerate
    generate 
        localparam integer d193 = 25;
        for (n193 = 0; n193 < 16; n193 = n193 + 1) 
        begin: outbit193
            assign data_11[n193 + d193*16 + c6*28*16] = data_11_array[c6][d193][n193];
        end
    endgenerate
    generate 
        localparam integer d194 = 26;
        for (n194 = 0; n194 < 16; n194 = n194 + 1) 
        begin: outbit194
            assign data_11[n194 + d194*16 + c6*28*16] = data_11_array[c6][d194][n194];
        end
    endgenerate
    generate 
        localparam integer d195 = 27;
        for (n195 = 0; n195 < 16; n195 = n195 + 1) 
        begin: outbit195
            assign data_11[n195 + d195*16 + c6*28*16] = data_11_array[c6][d195][n195];
        end
    endgenerate
    localparam integer c7 = 7;
    generate 
        localparam integer d196 = 0;
        for (n196 = 0; n196 < 16; n196 = n196 + 1) 
        begin: outbit196
            assign data_11[n196 + d196*16 + c7*28*16] = data_11_array[c7][d196][n196];
        end
    endgenerate
    generate 
        localparam integer d197 = 1;
        for (n197 = 0; n197 < 16; n197 = n197 + 1) 
        begin: outbit197
            assign data_11[n197 + d197*16 + c7*28*16] = data_11_array[c7][d197][n197];
        end
    endgenerate
    generate 
        localparam integer d198 = 2;
        for (n198 = 0; n198 < 16; n198 = n198 + 1) 
        begin: outbit198
            assign data_11[n198 + d198*16 + c7*28*16] = data_11_array[c7][d198][n198];
        end
    endgenerate
    generate 
        localparam integer d199 = 3;
        for (n199 = 0; n199 < 16; n199 = n199 + 1) 
        begin: outbit199
            assign data_11[n199 + d199*16 + c7*28*16] = data_11_array[c7][d199][n199];
        end
    endgenerate
    generate 
        localparam integer d200 = 4;
        for (n200 = 0; n200 < 16; n200 = n200 + 1) 
        begin: outbit200
            assign data_11[n200 + d200*16 + c7*28*16] = data_11_array[c7][d200][n200];
        end
    endgenerate
    generate 
        localparam integer d201 = 5;
        for (n201 = 0; n201 < 16; n201 = n201 + 1) 
        begin: outbit201
            assign data_11[n201 + d201*16 + c7*28*16] = data_11_array[c7][d201][n201];
        end
    endgenerate
    generate 
        localparam integer d202 = 6;
        for (n202 = 0; n202 < 16; n202 = n202 + 1) 
        begin: outbit202
            assign data_11[n202 + d202*16 + c7*28*16] = data_11_array[c7][d202][n202];
        end
    endgenerate
    generate 
        localparam integer d203 = 7;
        for (n203 = 0; n203 < 16; n203 = n203 + 1) 
        begin: outbit203
            assign data_11[n203 + d203*16 + c7*28*16] = data_11_array[c7][d203][n203];
        end
    endgenerate
    generate 
        localparam integer d204 = 8;
        for (n204 = 0; n204 < 16; n204 = n204 + 1) 
        begin: outbit204
            assign data_11[n204 + d204*16 + c7*28*16] = data_11_array[c7][d204][n204];
        end
    endgenerate
    generate 
        localparam integer d205 = 9;
        for (n205 = 0; n205 < 16; n205 = n205 + 1) 
        begin: outbit205
            assign data_11[n205 + d205*16 + c7*28*16] = data_11_array[c7][d205][n205];
        end
    endgenerate
    generate 
        localparam integer d206 = 10;
        for (n206 = 0; n206 < 16; n206 = n206 + 1) 
        begin: outbit206
            assign data_11[n206 + d206*16 + c7*28*16] = data_11_array[c7][d206][n206];
        end
    endgenerate
    generate 
        localparam integer d207 = 11;
        for (n207 = 0; n207 < 16; n207 = n207 + 1) 
        begin: outbit207
            assign data_11[n207 + d207*16 + c7*28*16] = data_11_array[c7][d207][n207];
        end
    endgenerate
    generate 
        localparam integer d208 = 12;
        for (n208 = 0; n208 < 16; n208 = n208 + 1) 
        begin: outbit208
            assign data_11[n208 + d208*16 + c7*28*16] = data_11_array[c7][d208][n208];
        end
    endgenerate
    generate 
        localparam integer d209 = 13;
        for (n209 = 0; n209 < 16; n209 = n209 + 1) 
        begin: outbit209
            assign data_11[n209 + d209*16 + c7*28*16] = data_11_array[c7][d209][n209];
        end
    endgenerate
    generate 
        localparam integer d210 = 14;
        for (n210 = 0; n210 < 16; n210 = n210 + 1) 
        begin: outbit210
            assign data_11[n210 + d210*16 + c7*28*16] = data_11_array[c7][d210][n210];
        end
    endgenerate
    generate 
        localparam integer d211 = 15;
        for (n211 = 0; n211 < 16; n211 = n211 + 1) 
        begin: outbit211
            assign data_11[n211 + d211*16 + c7*28*16] = data_11_array[c7][d211][n211];
        end
    endgenerate
    generate 
        localparam integer d212 = 16;
        for (n212 = 0; n212 < 16; n212 = n212 + 1) 
        begin: outbit212
            assign data_11[n212 + d212*16 + c7*28*16] = data_11_array[c7][d212][n212];
        end
    endgenerate
    generate 
        localparam integer d213 = 17;
        for (n213 = 0; n213 < 16; n213 = n213 + 1) 
        begin: outbit213
            assign data_11[n213 + d213*16 + c7*28*16] = data_11_array[c7][d213][n213];
        end
    endgenerate
    generate 
        localparam integer d214 = 18;
        for (n214 = 0; n214 < 16; n214 = n214 + 1) 
        begin: outbit214
            assign data_11[n214 + d214*16 + c7*28*16] = data_11_array[c7][d214][n214];
        end
    endgenerate
    generate 
        localparam integer d215 = 19;
        for (n215 = 0; n215 < 16; n215 = n215 + 1) 
        begin: outbit215
            assign data_11[n215 + d215*16 + c7*28*16] = data_11_array[c7][d215][n215];
        end
    endgenerate
    generate 
        localparam integer d216 = 20;
        for (n216 = 0; n216 < 16; n216 = n216 + 1) 
        begin: outbit216
            assign data_11[n216 + d216*16 + c7*28*16] = data_11_array[c7][d216][n216];
        end
    endgenerate
    generate 
        localparam integer d217 = 21;
        for (n217 = 0; n217 < 16; n217 = n217 + 1) 
        begin: outbit217
            assign data_11[n217 + d217*16 + c7*28*16] = data_11_array[c7][d217][n217];
        end
    endgenerate
    generate 
        localparam integer d218 = 22;
        for (n218 = 0; n218 < 16; n218 = n218 + 1) 
        begin: outbit218
            assign data_11[n218 + d218*16 + c7*28*16] = data_11_array[c7][d218][n218];
        end
    endgenerate
    generate 
        localparam integer d219 = 23;
        for (n219 = 0; n219 < 16; n219 = n219 + 1) 
        begin: outbit219
            assign data_11[n219 + d219*16 + c7*28*16] = data_11_array[c7][d219][n219];
        end
    endgenerate
    generate 
        localparam integer d220 = 24;
        for (n220 = 0; n220 < 16; n220 = n220 + 1) 
        begin: outbit220
            assign data_11[n220 + d220*16 + c7*28*16] = data_11_array[c7][d220][n220];
        end
    endgenerate
    generate 
        localparam integer d221 = 25;
        for (n221 = 0; n221 < 16; n221 = n221 + 1) 
        begin: outbit221
            assign data_11[n221 + d221*16 + c7*28*16] = data_11_array[c7][d221][n221];
        end
    endgenerate
    generate 
        localparam integer d222 = 26;
        for (n222 = 0; n222 < 16; n222 = n222 + 1) 
        begin: outbit222
            assign data_11[n222 + d222*16 + c7*28*16] = data_11_array[c7][d222][n222];
        end
    endgenerate
    generate 
        localparam integer d223 = 27;
        for (n223 = 0; n223 < 16; n223 = n223 + 1) 
        begin: outbit223
            assign data_11[n223 + d223*16 + c7*28*16] = data_11_array[c7][d223][n223];
        end
    endgenerate
    localparam integer c8 = 8;
    generate 
        localparam integer d224 = 0;
        for (n224 = 0; n224 < 16; n224 = n224 + 1) 
        begin: outbit224
            assign data_11[n224 + d224*16 + c8*28*16] = data_11_array[c8][d224][n224];
        end
    endgenerate
    generate 
        localparam integer d225 = 1;
        for (n225 = 0; n225 < 16; n225 = n225 + 1) 
        begin: outbit225
            assign data_11[n225 + d225*16 + c8*28*16] = data_11_array[c8][d225][n225];
        end
    endgenerate
    generate 
        localparam integer d226 = 2;
        for (n226 = 0; n226 < 16; n226 = n226 + 1) 
        begin: outbit226
            assign data_11[n226 + d226*16 + c8*28*16] = data_11_array[c8][d226][n226];
        end
    endgenerate
    generate 
        localparam integer d227 = 3;
        for (n227 = 0; n227 < 16; n227 = n227 + 1) 
        begin: outbit227
            assign data_11[n227 + d227*16 + c8*28*16] = data_11_array[c8][d227][n227];
        end
    endgenerate
    generate 
        localparam integer d228 = 4;
        for (n228 = 0; n228 < 16; n228 = n228 + 1) 
        begin: outbit228
            assign data_11[n228 + d228*16 + c8*28*16] = data_11_array[c8][d228][n228];
        end
    endgenerate
    generate 
        localparam integer d229 = 5;
        for (n229 = 0; n229 < 16; n229 = n229 + 1) 
        begin: outbit229
            assign data_11[n229 + d229*16 + c8*28*16] = data_11_array[c8][d229][n229];
        end
    endgenerate
    generate 
        localparam integer d230 = 6;
        for (n230 = 0; n230 < 16; n230 = n230 + 1) 
        begin: outbit230
            assign data_11[n230 + d230*16 + c8*28*16] = data_11_array[c8][d230][n230];
        end
    endgenerate
    generate 
        localparam integer d231 = 7;
        for (n231 = 0; n231 < 16; n231 = n231 + 1) 
        begin: outbit231
            assign data_11[n231 + d231*16 + c8*28*16] = data_11_array[c8][d231][n231];
        end
    endgenerate
    generate 
        localparam integer d232 = 8;
        for (n232 = 0; n232 < 16; n232 = n232 + 1) 
        begin: outbit232
            assign data_11[n232 + d232*16 + c8*28*16] = data_11_array[c8][d232][n232];
        end
    endgenerate
    generate 
        localparam integer d233 = 9;
        for (n233 = 0; n233 < 16; n233 = n233 + 1) 
        begin: outbit233
            assign data_11[n233 + d233*16 + c8*28*16] = data_11_array[c8][d233][n233];
        end
    endgenerate
    generate 
        localparam integer d234 = 10;
        for (n234 = 0; n234 < 16; n234 = n234 + 1) 
        begin: outbit234
            assign data_11[n234 + d234*16 + c8*28*16] = data_11_array[c8][d234][n234];
        end
    endgenerate
    generate 
        localparam integer d235 = 11;
        for (n235 = 0; n235 < 16; n235 = n235 + 1) 
        begin: outbit235
            assign data_11[n235 + d235*16 + c8*28*16] = data_11_array[c8][d235][n235];
        end
    endgenerate
    generate 
        localparam integer d236 = 12;
        for (n236 = 0; n236 < 16; n236 = n236 + 1) 
        begin: outbit236
            assign data_11[n236 + d236*16 + c8*28*16] = data_11_array[c8][d236][n236];
        end
    endgenerate
    generate 
        localparam integer d237 = 13;
        for (n237 = 0; n237 < 16; n237 = n237 + 1) 
        begin: outbit237
            assign data_11[n237 + d237*16 + c8*28*16] = data_11_array[c8][d237][n237];
        end
    endgenerate
    generate 
        localparam integer d238 = 14;
        for (n238 = 0; n238 < 16; n238 = n238 + 1) 
        begin: outbit238
            assign data_11[n238 + d238*16 + c8*28*16] = data_11_array[c8][d238][n238];
        end
    endgenerate
    generate 
        localparam integer d239 = 15;
        for (n239 = 0; n239 < 16; n239 = n239 + 1) 
        begin: outbit239
            assign data_11[n239 + d239*16 + c8*28*16] = data_11_array[c8][d239][n239];
        end
    endgenerate
    generate 
        localparam integer d240 = 16;
        for (n240 = 0; n240 < 16; n240 = n240 + 1) 
        begin: outbit240
            assign data_11[n240 + d240*16 + c8*28*16] = data_11_array[c8][d240][n240];
        end
    endgenerate
    generate 
        localparam integer d241 = 17;
        for (n241 = 0; n241 < 16; n241 = n241 + 1) 
        begin: outbit241
            assign data_11[n241 + d241*16 + c8*28*16] = data_11_array[c8][d241][n241];
        end
    endgenerate
    generate 
        localparam integer d242 = 18;
        for (n242 = 0; n242 < 16; n242 = n242 + 1) 
        begin: outbit242
            assign data_11[n242 + d242*16 + c8*28*16] = data_11_array[c8][d242][n242];
        end
    endgenerate
    generate 
        localparam integer d243 = 19;
        for (n243 = 0; n243 < 16; n243 = n243 + 1) 
        begin: outbit243
            assign data_11[n243 + d243*16 + c8*28*16] = data_11_array[c8][d243][n243];
        end
    endgenerate
    generate 
        localparam integer d244 = 20;
        for (n244 = 0; n244 < 16; n244 = n244 + 1) 
        begin: outbit244
            assign data_11[n244 + d244*16 + c8*28*16] = data_11_array[c8][d244][n244];
        end
    endgenerate
    generate 
        localparam integer d245 = 21;
        for (n245 = 0; n245 < 16; n245 = n245 + 1) 
        begin: outbit245
            assign data_11[n245 + d245*16 + c8*28*16] = data_11_array[c8][d245][n245];
        end
    endgenerate
    generate 
        localparam integer d246 = 22;
        for (n246 = 0; n246 < 16; n246 = n246 + 1) 
        begin: outbit246
            assign data_11[n246 + d246*16 + c8*28*16] = data_11_array[c8][d246][n246];
        end
    endgenerate
    generate 
        localparam integer d247 = 23;
        for (n247 = 0; n247 < 16; n247 = n247 + 1) 
        begin: outbit247
            assign data_11[n247 + d247*16 + c8*28*16] = data_11_array[c8][d247][n247];
        end
    endgenerate
    generate 
        localparam integer d248 = 24;
        for (n248 = 0; n248 < 16; n248 = n248 + 1) 
        begin: outbit248
            assign data_11[n248 + d248*16 + c8*28*16] = data_11_array[c8][d248][n248];
        end
    endgenerate
    generate 
        localparam integer d249 = 25;
        for (n249 = 0; n249 < 16; n249 = n249 + 1) 
        begin: outbit249
            assign data_11[n249 + d249*16 + c8*28*16] = data_11_array[c8][d249][n249];
        end
    endgenerate
    generate 
        localparam integer d250 = 26;
        for (n250 = 0; n250 < 16; n250 = n250 + 1) 
        begin: outbit250
            assign data_11[n250 + d250*16 + c8*28*16] = data_11_array[c8][d250][n250];
        end
    endgenerate
    generate 
        localparam integer d251 = 27;
        for (n251 = 0; n251 < 16; n251 = n251 + 1) 
        begin: outbit251
            assign data_11[n251 + d251*16 + c8*28*16] = data_11_array[c8][d251][n251];
        end
    endgenerate
    localparam integer c9 = 9;
    generate 
        localparam integer d252 = 0;
        for (n252 = 0; n252 < 16; n252 = n252 + 1) 
        begin: outbit252
            assign data_11[n252 + d252*16 + c9*28*16] = data_11_array[c9][d252][n252];
        end
    endgenerate
    generate 
        localparam integer d253 = 1;
        for (n253 = 0; n253 < 16; n253 = n253 + 1) 
        begin: outbit253
            assign data_11[n253 + d253*16 + c9*28*16] = data_11_array[c9][d253][n253];
        end
    endgenerate
    generate 
        localparam integer d254 = 2;
        for (n254 = 0; n254 < 16; n254 = n254 + 1) 
        begin: outbit254
            assign data_11[n254 + d254*16 + c9*28*16] = data_11_array[c9][d254][n254];
        end
    endgenerate
    generate 
        localparam integer d255 = 3;
        for (n255 = 0; n255 < 16; n255 = n255 + 1) 
        begin: outbit255
            assign data_11[n255 + d255*16 + c9*28*16] = data_11_array[c9][d255][n255];
        end
    endgenerate
    generate 
        localparam integer d256 = 4;
        for (n256 = 0; n256 < 16; n256 = n256 + 1) 
        begin: outbit256
            assign data_11[n256 + d256*16 + c9*28*16] = data_11_array[c9][d256][n256];
        end
    endgenerate
    generate 
        localparam integer d257 = 5;
        for (n257 = 0; n257 < 16; n257 = n257 + 1) 
        begin: outbit257
            assign data_11[n257 + d257*16 + c9*28*16] = data_11_array[c9][d257][n257];
        end
    endgenerate
    generate 
        localparam integer d258 = 6;
        for (n258 = 0; n258 < 16; n258 = n258 + 1) 
        begin: outbit258
            assign data_11[n258 + d258*16 + c9*28*16] = data_11_array[c9][d258][n258];
        end
    endgenerate
    generate 
        localparam integer d259 = 7;
        for (n259 = 0; n259 < 16; n259 = n259 + 1) 
        begin: outbit259
            assign data_11[n259 + d259*16 + c9*28*16] = data_11_array[c9][d259][n259];
        end
    endgenerate
    generate 
        localparam integer d260 = 8;
        for (n260 = 0; n260 < 16; n260 = n260 + 1) 
        begin: outbit260
            assign data_11[n260 + d260*16 + c9*28*16] = data_11_array[c9][d260][n260];
        end
    endgenerate
    generate 
        localparam integer d261 = 9;
        for (n261 = 0; n261 < 16; n261 = n261 + 1) 
        begin: outbit261
            assign data_11[n261 + d261*16 + c9*28*16] = data_11_array[c9][d261][n261];
        end
    endgenerate
    generate 
        localparam integer d262 = 10;
        for (n262 = 0; n262 < 16; n262 = n262 + 1) 
        begin: outbit262
            assign data_11[n262 + d262*16 + c9*28*16] = data_11_array[c9][d262][n262];
        end
    endgenerate
    generate 
        localparam integer d263 = 11;
        for (n263 = 0; n263 < 16; n263 = n263 + 1) 
        begin: outbit263
            assign data_11[n263 + d263*16 + c9*28*16] = data_11_array[c9][d263][n263];
        end
    endgenerate
    generate 
        localparam integer d264 = 12;
        for (n264 = 0; n264 < 16; n264 = n264 + 1) 
        begin: outbit264
            assign data_11[n264 + d264*16 + c9*28*16] = data_11_array[c9][d264][n264];
        end
    endgenerate
    generate 
        localparam integer d265 = 13;
        for (n265 = 0; n265 < 16; n265 = n265 + 1) 
        begin: outbit265
            assign data_11[n265 + d265*16 + c9*28*16] = data_11_array[c9][d265][n265];
        end
    endgenerate
    generate 
        localparam integer d266 = 14;
        for (n266 = 0; n266 < 16; n266 = n266 + 1) 
        begin: outbit266
            assign data_11[n266 + d266*16 + c9*28*16] = data_11_array[c9][d266][n266];
        end
    endgenerate
    generate 
        localparam integer d267 = 15;
        for (n267 = 0; n267 < 16; n267 = n267 + 1) 
        begin: outbit267
            assign data_11[n267 + d267*16 + c9*28*16] = data_11_array[c9][d267][n267];
        end
    endgenerate
    generate 
        localparam integer d268 = 16;
        for (n268 = 0; n268 < 16; n268 = n268 + 1) 
        begin: outbit268
            assign data_11[n268 + d268*16 + c9*28*16] = data_11_array[c9][d268][n268];
        end
    endgenerate
    generate 
        localparam integer d269 = 17;
        for (n269 = 0; n269 < 16; n269 = n269 + 1) 
        begin: outbit269
            assign data_11[n269 + d269*16 + c9*28*16] = data_11_array[c9][d269][n269];
        end
    endgenerate
    generate 
        localparam integer d270 = 18;
        for (n270 = 0; n270 < 16; n270 = n270 + 1) 
        begin: outbit270
            assign data_11[n270 + d270*16 + c9*28*16] = data_11_array[c9][d270][n270];
        end
    endgenerate
    generate 
        localparam integer d271 = 19;
        for (n271 = 0; n271 < 16; n271 = n271 + 1) 
        begin: outbit271
            assign data_11[n271 + d271*16 + c9*28*16] = data_11_array[c9][d271][n271];
        end
    endgenerate
    generate 
        localparam integer d272 = 20;
        for (n272 = 0; n272 < 16; n272 = n272 + 1) 
        begin: outbit272
            assign data_11[n272 + d272*16 + c9*28*16] = data_11_array[c9][d272][n272];
        end
    endgenerate
    generate 
        localparam integer d273 = 21;
        for (n273 = 0; n273 < 16; n273 = n273 + 1) 
        begin: outbit273
            assign data_11[n273 + d273*16 + c9*28*16] = data_11_array[c9][d273][n273];
        end
    endgenerate
    generate 
        localparam integer d274 = 22;
        for (n274 = 0; n274 < 16; n274 = n274 + 1) 
        begin: outbit274
            assign data_11[n274 + d274*16 + c9*28*16] = data_11_array[c9][d274][n274];
        end
    endgenerate
    generate 
        localparam integer d275 = 23;
        for (n275 = 0; n275 < 16; n275 = n275 + 1) 
        begin: outbit275
            assign data_11[n275 + d275*16 + c9*28*16] = data_11_array[c9][d275][n275];
        end
    endgenerate
    generate 
        localparam integer d276 = 24;
        for (n276 = 0; n276 < 16; n276 = n276 + 1) 
        begin: outbit276
            assign data_11[n276 + d276*16 + c9*28*16] = data_11_array[c9][d276][n276];
        end
    endgenerate
    generate 
        localparam integer d277 = 25;
        for (n277 = 0; n277 < 16; n277 = n277 + 1) 
        begin: outbit277
            assign data_11[n277 + d277*16 + c9*28*16] = data_11_array[c9][d277][n277];
        end
    endgenerate
    generate 
        localparam integer d278 = 26;
        for (n278 = 0; n278 < 16; n278 = n278 + 1) 
        begin: outbit278
            assign data_11[n278 + d278*16 + c9*28*16] = data_11_array[c9][d278][n278];
        end
    endgenerate
    generate 
        localparam integer d279 = 27;
        for (n279 = 0; n279 < 16; n279 = n279 + 1) 
        begin: outbit279
            assign data_11[n279 + d279*16 + c9*28*16] = data_11_array[c9][d279][n279];
        end
    endgenerate
    localparam integer c10 = 10;
    generate 
        localparam integer d280 = 0;
        for (n280 = 0; n280 < 16; n280 = n280 + 1) 
        begin: outbit280
            assign data_11[n280 + d280*16 + c10*28*16] = data_11_array[c10][d280][n280];
        end
    endgenerate
    generate 
        localparam integer d281 = 1;
        for (n281 = 0; n281 < 16; n281 = n281 + 1) 
        begin: outbit281
            assign data_11[n281 + d281*16 + c10*28*16] = data_11_array[c10][d281][n281];
        end
    endgenerate
    generate 
        localparam integer d282 = 2;
        for (n282 = 0; n282 < 16; n282 = n282 + 1) 
        begin: outbit282
            assign data_11[n282 + d282*16 + c10*28*16] = data_11_array[c10][d282][n282];
        end
    endgenerate
    generate 
        localparam integer d283 = 3;
        for (n283 = 0; n283 < 16; n283 = n283 + 1) 
        begin: outbit283
            assign data_11[n283 + d283*16 + c10*28*16] = data_11_array[c10][d283][n283];
        end
    endgenerate
    generate 
        localparam integer d284 = 4;
        for (n284 = 0; n284 < 16; n284 = n284 + 1) 
        begin: outbit284
            assign data_11[n284 + d284*16 + c10*28*16] = data_11_array[c10][d284][n284];
        end
    endgenerate
    generate 
        localparam integer d285 = 5;
        for (n285 = 0; n285 < 16; n285 = n285 + 1) 
        begin: outbit285
            assign data_11[n285 + d285*16 + c10*28*16] = data_11_array[c10][d285][n285];
        end
    endgenerate
    generate 
        localparam integer d286 = 6;
        for (n286 = 0; n286 < 16; n286 = n286 + 1) 
        begin: outbit286
            assign data_11[n286 + d286*16 + c10*28*16] = data_11_array[c10][d286][n286];
        end
    endgenerate
    generate 
        localparam integer d287 = 7;
        for (n287 = 0; n287 < 16; n287 = n287 + 1) 
        begin: outbit287
            assign data_11[n287 + d287*16 + c10*28*16] = data_11_array[c10][d287][n287];
        end
    endgenerate
    generate 
        localparam integer d288 = 8;
        for (n288 = 0; n288 < 16; n288 = n288 + 1) 
        begin: outbit288
            assign data_11[n288 + d288*16 + c10*28*16] = data_11_array[c10][d288][n288];
        end
    endgenerate
    generate 
        localparam integer d289 = 9;
        for (n289 = 0; n289 < 16; n289 = n289 + 1) 
        begin: outbit289
            assign data_11[n289 + d289*16 + c10*28*16] = data_11_array[c10][d289][n289];
        end
    endgenerate
    generate 
        localparam integer d290 = 10;
        for (n290 = 0; n290 < 16; n290 = n290 + 1) 
        begin: outbit290
            assign data_11[n290 + d290*16 + c10*28*16] = data_11_array[c10][d290][n290];
        end
    endgenerate
    generate 
        localparam integer d291 = 11;
        for (n291 = 0; n291 < 16; n291 = n291 + 1) 
        begin: outbit291
            assign data_11[n291 + d291*16 + c10*28*16] = data_11_array[c10][d291][n291];
        end
    endgenerate
    generate 
        localparam integer d292 = 12;
        for (n292 = 0; n292 < 16; n292 = n292 + 1) 
        begin: outbit292
            assign data_11[n292 + d292*16 + c10*28*16] = data_11_array[c10][d292][n292];
        end
    endgenerate
    generate 
        localparam integer d293 = 13;
        for (n293 = 0; n293 < 16; n293 = n293 + 1) 
        begin: outbit293
            assign data_11[n293 + d293*16 + c10*28*16] = data_11_array[c10][d293][n293];
        end
    endgenerate
    generate 
        localparam integer d294 = 14;
        for (n294 = 0; n294 < 16; n294 = n294 + 1) 
        begin: outbit294
            assign data_11[n294 + d294*16 + c10*28*16] = data_11_array[c10][d294][n294];
        end
    endgenerate
    generate 
        localparam integer d295 = 15;
        for (n295 = 0; n295 < 16; n295 = n295 + 1) 
        begin: outbit295
            assign data_11[n295 + d295*16 + c10*28*16] = data_11_array[c10][d295][n295];
        end
    endgenerate
    generate 
        localparam integer d296 = 16;
        for (n296 = 0; n296 < 16; n296 = n296 + 1) 
        begin: outbit296
            assign data_11[n296 + d296*16 + c10*28*16] = data_11_array[c10][d296][n296];
        end
    endgenerate
    generate 
        localparam integer d297 = 17;
        for (n297 = 0; n297 < 16; n297 = n297 + 1) 
        begin: outbit297
            assign data_11[n297 + d297*16 + c10*28*16] = data_11_array[c10][d297][n297];
        end
    endgenerate
    generate 
        localparam integer d298 = 18;
        for (n298 = 0; n298 < 16; n298 = n298 + 1) 
        begin: outbit298
            assign data_11[n298 + d298*16 + c10*28*16] = data_11_array[c10][d298][n298];
        end
    endgenerate
    generate 
        localparam integer d299 = 19;
        for (n299 = 0; n299 < 16; n299 = n299 + 1) 
        begin: outbit299
            assign data_11[n299 + d299*16 + c10*28*16] = data_11_array[c10][d299][n299];
        end
    endgenerate
    generate 
        localparam integer d300 = 20;
        for (n300 = 0; n300 < 16; n300 = n300 + 1) 
        begin: outbit300
            assign data_11[n300 + d300*16 + c10*28*16] = data_11_array[c10][d300][n300];
        end
    endgenerate
    generate 
        localparam integer d301 = 21;
        for (n301 = 0; n301 < 16; n301 = n301 + 1) 
        begin: outbit301
            assign data_11[n301 + d301*16 + c10*28*16] = data_11_array[c10][d301][n301];
        end
    endgenerate
    generate 
        localparam integer d302 = 22;
        for (n302 = 0; n302 < 16; n302 = n302 + 1) 
        begin: outbit302
            assign data_11[n302 + d302*16 + c10*28*16] = data_11_array[c10][d302][n302];
        end
    endgenerate
    generate 
        localparam integer d303 = 23;
        for (n303 = 0; n303 < 16; n303 = n303 + 1) 
        begin: outbit303
            assign data_11[n303 + d303*16 + c10*28*16] = data_11_array[c10][d303][n303];
        end
    endgenerate
    generate 
        localparam integer d304 = 24;
        for (n304 = 0; n304 < 16; n304 = n304 + 1) 
        begin: outbit304
            assign data_11[n304 + d304*16 + c10*28*16] = data_11_array[c10][d304][n304];
        end
    endgenerate
    generate 
        localparam integer d305 = 25;
        for (n305 = 0; n305 < 16; n305 = n305 + 1) 
        begin: outbit305
            assign data_11[n305 + d305*16 + c10*28*16] = data_11_array[c10][d305][n305];
        end
    endgenerate
    generate 
        localparam integer d306 = 26;
        for (n306 = 0; n306 < 16; n306 = n306 + 1) 
        begin: outbit306
            assign data_11[n306 + d306*16 + c10*28*16] = data_11_array[c10][d306][n306];
        end
    endgenerate
    generate 
        localparam integer d307 = 27;
        for (n307 = 0; n307 < 16; n307 = n307 + 1) 
        begin: outbit307
            assign data_11[n307 + d307*16 + c10*28*16] = data_11_array[c10][d307][n307];
        end
    endgenerate
    localparam integer c11 = 11;
    generate 
        localparam integer d308 = 0;
        for (n308 = 0; n308 < 16; n308 = n308 + 1) 
        begin: outbit308
            assign data_11[n308 + d308*16 + c11*28*16] = data_11_array[c11][d308][n308];
        end
    endgenerate
    generate 
        localparam integer d309 = 1;
        for (n309 = 0; n309 < 16; n309 = n309 + 1) 
        begin: outbit309
            assign data_11[n309 + d309*16 + c11*28*16] = data_11_array[c11][d309][n309];
        end
    endgenerate
    generate 
        localparam integer d310 = 2;
        for (n310 = 0; n310 < 16; n310 = n310 + 1) 
        begin: outbit310
            assign data_11[n310 + d310*16 + c11*28*16] = data_11_array[c11][d310][n310];
        end
    endgenerate
    generate 
        localparam integer d311 = 3;
        for (n311 = 0; n311 < 16; n311 = n311 + 1) 
        begin: outbit311
            assign data_11[n311 + d311*16 + c11*28*16] = data_11_array[c11][d311][n311];
        end
    endgenerate
    generate 
        localparam integer d312 = 4;
        for (n312 = 0; n312 < 16; n312 = n312 + 1) 
        begin: outbit312
            assign data_11[n312 + d312*16 + c11*28*16] = data_11_array[c11][d312][n312];
        end
    endgenerate
    generate 
        localparam integer d313 = 5;
        for (n313 = 0; n313 < 16; n313 = n313 + 1) 
        begin: outbit313
            assign data_11[n313 + d313*16 + c11*28*16] = data_11_array[c11][d313][n313];
        end
    endgenerate
    generate 
        localparam integer d314 = 6;
        for (n314 = 0; n314 < 16; n314 = n314 + 1) 
        begin: outbit314
            assign data_11[n314 + d314*16 + c11*28*16] = data_11_array[c11][d314][n314];
        end
    endgenerate
    generate 
        localparam integer d315 = 7;
        for (n315 = 0; n315 < 16; n315 = n315 + 1) 
        begin: outbit315
            assign data_11[n315 + d315*16 + c11*28*16] = data_11_array[c11][d315][n315];
        end
    endgenerate
    generate 
        localparam integer d316 = 8;
        for (n316 = 0; n316 < 16; n316 = n316 + 1) 
        begin: outbit316
            assign data_11[n316 + d316*16 + c11*28*16] = data_11_array[c11][d316][n316];
        end
    endgenerate
    generate 
        localparam integer d317 = 9;
        for (n317 = 0; n317 < 16; n317 = n317 + 1) 
        begin: outbit317
            assign data_11[n317 + d317*16 + c11*28*16] = data_11_array[c11][d317][n317];
        end
    endgenerate
    generate 
        localparam integer d318 = 10;
        for (n318 = 0; n318 < 16; n318 = n318 + 1) 
        begin: outbit318
            assign data_11[n318 + d318*16 + c11*28*16] = data_11_array[c11][d318][n318];
        end
    endgenerate
    generate 
        localparam integer d319 = 11;
        for (n319 = 0; n319 < 16; n319 = n319 + 1) 
        begin: outbit319
            assign data_11[n319 + d319*16 + c11*28*16] = data_11_array[c11][d319][n319];
        end
    endgenerate
    generate 
        localparam integer d320 = 12;
        for (n320 = 0; n320 < 16; n320 = n320 + 1) 
        begin: outbit320
            assign data_11[n320 + d320*16 + c11*28*16] = data_11_array[c11][d320][n320];
        end
    endgenerate
    generate 
        localparam integer d321 = 13;
        for (n321 = 0; n321 < 16; n321 = n321 + 1) 
        begin: outbit321
            assign data_11[n321 + d321*16 + c11*28*16] = data_11_array[c11][d321][n321];
        end
    endgenerate
    generate 
        localparam integer d322 = 14;
        for (n322 = 0; n322 < 16; n322 = n322 + 1) 
        begin: outbit322
            assign data_11[n322 + d322*16 + c11*28*16] = data_11_array[c11][d322][n322];
        end
    endgenerate
    generate 
        localparam integer d323 = 15;
        for (n323 = 0; n323 < 16; n323 = n323 + 1) 
        begin: outbit323
            assign data_11[n323 + d323*16 + c11*28*16] = data_11_array[c11][d323][n323];
        end
    endgenerate
    generate 
        localparam integer d324 = 16;
        for (n324 = 0; n324 < 16; n324 = n324 + 1) 
        begin: outbit324
            assign data_11[n324 + d324*16 + c11*28*16] = data_11_array[c11][d324][n324];
        end
    endgenerate
    generate 
        localparam integer d325 = 17;
        for (n325 = 0; n325 < 16; n325 = n325 + 1) 
        begin: outbit325
            assign data_11[n325 + d325*16 + c11*28*16] = data_11_array[c11][d325][n325];
        end
    endgenerate
    generate 
        localparam integer d326 = 18;
        for (n326 = 0; n326 < 16; n326 = n326 + 1) 
        begin: outbit326
            assign data_11[n326 + d326*16 + c11*28*16] = data_11_array[c11][d326][n326];
        end
    endgenerate
    generate 
        localparam integer d327 = 19;
        for (n327 = 0; n327 < 16; n327 = n327 + 1) 
        begin: outbit327
            assign data_11[n327 + d327*16 + c11*28*16] = data_11_array[c11][d327][n327];
        end
    endgenerate
    generate 
        localparam integer d328 = 20;
        for (n328 = 0; n328 < 16; n328 = n328 + 1) 
        begin: outbit328
            assign data_11[n328 + d328*16 + c11*28*16] = data_11_array[c11][d328][n328];
        end
    endgenerate
    generate 
        localparam integer d329 = 21;
        for (n329 = 0; n329 < 16; n329 = n329 + 1) 
        begin: outbit329
            assign data_11[n329 + d329*16 + c11*28*16] = data_11_array[c11][d329][n329];
        end
    endgenerate
    generate 
        localparam integer d330 = 22;
        for (n330 = 0; n330 < 16; n330 = n330 + 1) 
        begin: outbit330
            assign data_11[n330 + d330*16 + c11*28*16] = data_11_array[c11][d330][n330];
        end
    endgenerate
    generate 
        localparam integer d331 = 23;
        for (n331 = 0; n331 < 16; n331 = n331 + 1) 
        begin: outbit331
            assign data_11[n331 + d331*16 + c11*28*16] = data_11_array[c11][d331][n331];
        end
    endgenerate
    generate 
        localparam integer d332 = 24;
        for (n332 = 0; n332 < 16; n332 = n332 + 1) 
        begin: outbit332
            assign data_11[n332 + d332*16 + c11*28*16] = data_11_array[c11][d332][n332];
        end
    endgenerate
    generate 
        localparam integer d333 = 25;
        for (n333 = 0; n333 < 16; n333 = n333 + 1) 
        begin: outbit333
            assign data_11[n333 + d333*16 + c11*28*16] = data_11_array[c11][d333][n333];
        end
    endgenerate
    generate 
        localparam integer d334 = 26;
        for (n334 = 0; n334 < 16; n334 = n334 + 1) 
        begin: outbit334
            assign data_11[n334 + d334*16 + c11*28*16] = data_11_array[c11][d334][n334];
        end
    endgenerate
    generate 
        localparam integer d335 = 27;
        for (n335 = 0; n335 < 16; n335 = n335 + 1) 
        begin: outbit335
            assign data_11[n335 + d335*16 + c11*28*16] = data_11_array[c11][d335][n335];
        end
    endgenerate
    localparam integer c12 = 12;
    generate 
        localparam integer d336 = 0;
        for (n336 = 0; n336 < 16; n336 = n336 + 1) 
        begin: outbit336
            assign data_11[n336 + d336*16 + c12*28*16] = data_11_array[c12][d336][n336];
        end
    endgenerate
    generate 
        localparam integer d337 = 1;
        for (n337 = 0; n337 < 16; n337 = n337 + 1) 
        begin: outbit337
            assign data_11[n337 + d337*16 + c12*28*16] = data_11_array[c12][d337][n337];
        end
    endgenerate
    generate 
        localparam integer d338 = 2;
        for (n338 = 0; n338 < 16; n338 = n338 + 1) 
        begin: outbit338
            assign data_11[n338 + d338*16 + c12*28*16] = data_11_array[c12][d338][n338];
        end
    endgenerate
    generate 
        localparam integer d339 = 3;
        for (n339 = 0; n339 < 16; n339 = n339 + 1) 
        begin: outbit339
            assign data_11[n339 + d339*16 + c12*28*16] = data_11_array[c12][d339][n339];
        end
    endgenerate
    generate 
        localparam integer d340 = 4;
        for (n340 = 0; n340 < 16; n340 = n340 + 1) 
        begin: outbit340
            assign data_11[n340 + d340*16 + c12*28*16] = data_11_array[c12][d340][n340];
        end
    endgenerate
    generate 
        localparam integer d341 = 5;
        for (n341 = 0; n341 < 16; n341 = n341 + 1) 
        begin: outbit341
            assign data_11[n341 + d341*16 + c12*28*16] = data_11_array[c12][d341][n341];
        end
    endgenerate
    generate 
        localparam integer d342 = 6;
        for (n342 = 0; n342 < 16; n342 = n342 + 1) 
        begin: outbit342
            assign data_11[n342 + d342*16 + c12*28*16] = data_11_array[c12][d342][n342];
        end
    endgenerate
    generate 
        localparam integer d343 = 7;
        for (n343 = 0; n343 < 16; n343 = n343 + 1) 
        begin: outbit343
            assign data_11[n343 + d343*16 + c12*28*16] = data_11_array[c12][d343][n343];
        end
    endgenerate
    generate 
        localparam integer d344 = 8;
        for (n344 = 0; n344 < 16; n344 = n344 + 1) 
        begin: outbit344
            assign data_11[n344 + d344*16 + c12*28*16] = data_11_array[c12][d344][n344];
        end
    endgenerate
    generate 
        localparam integer d345 = 9;
        for (n345 = 0; n345 < 16; n345 = n345 + 1) 
        begin: outbit345
            assign data_11[n345 + d345*16 + c12*28*16] = data_11_array[c12][d345][n345];
        end
    endgenerate
    generate 
        localparam integer d346 = 10;
        for (n346 = 0; n346 < 16; n346 = n346 + 1) 
        begin: outbit346
            assign data_11[n346 + d346*16 + c12*28*16] = data_11_array[c12][d346][n346];
        end
    endgenerate
    generate 
        localparam integer d347 = 11;
        for (n347 = 0; n347 < 16; n347 = n347 + 1) 
        begin: outbit347
            assign data_11[n347 + d347*16 + c12*28*16] = data_11_array[c12][d347][n347];
        end
    endgenerate
    generate 
        localparam integer d348 = 12;
        for (n348 = 0; n348 < 16; n348 = n348 + 1) 
        begin: outbit348
            assign data_11[n348 + d348*16 + c12*28*16] = data_11_array[c12][d348][n348];
        end
    endgenerate
    generate 
        localparam integer d349 = 13;
        for (n349 = 0; n349 < 16; n349 = n349 + 1) 
        begin: outbit349
            assign data_11[n349 + d349*16 + c12*28*16] = data_11_array[c12][d349][n349];
        end
    endgenerate
    generate 
        localparam integer d350 = 14;
        for (n350 = 0; n350 < 16; n350 = n350 + 1) 
        begin: outbit350
            assign data_11[n350 + d350*16 + c12*28*16] = data_11_array[c12][d350][n350];
        end
    endgenerate
    generate 
        localparam integer d351 = 15;
        for (n351 = 0; n351 < 16; n351 = n351 + 1) 
        begin: outbit351
            assign data_11[n351 + d351*16 + c12*28*16] = data_11_array[c12][d351][n351];
        end
    endgenerate
    generate 
        localparam integer d352 = 16;
        for (n352 = 0; n352 < 16; n352 = n352 + 1) 
        begin: outbit352
            assign data_11[n352 + d352*16 + c12*28*16] = data_11_array[c12][d352][n352];
        end
    endgenerate
    generate 
        localparam integer d353 = 17;
        for (n353 = 0; n353 < 16; n353 = n353 + 1) 
        begin: outbit353
            assign data_11[n353 + d353*16 + c12*28*16] = data_11_array[c12][d353][n353];
        end
    endgenerate
    generate 
        localparam integer d354 = 18;
        for (n354 = 0; n354 < 16; n354 = n354 + 1) 
        begin: outbit354
            assign data_11[n354 + d354*16 + c12*28*16] = data_11_array[c12][d354][n354];
        end
    endgenerate
    generate 
        localparam integer d355 = 19;
        for (n355 = 0; n355 < 16; n355 = n355 + 1) 
        begin: outbit355
            assign data_11[n355 + d355*16 + c12*28*16] = data_11_array[c12][d355][n355];
        end
    endgenerate
    generate 
        localparam integer d356 = 20;
        for (n356 = 0; n356 < 16; n356 = n356 + 1) 
        begin: outbit356
            assign data_11[n356 + d356*16 + c12*28*16] = data_11_array[c12][d356][n356];
        end
    endgenerate
    generate 
        localparam integer d357 = 21;
        for (n357 = 0; n357 < 16; n357 = n357 + 1) 
        begin: outbit357
            assign data_11[n357 + d357*16 + c12*28*16] = data_11_array[c12][d357][n357];
        end
    endgenerate
    generate 
        localparam integer d358 = 22;
        for (n358 = 0; n358 < 16; n358 = n358 + 1) 
        begin: outbit358
            assign data_11[n358 + d358*16 + c12*28*16] = data_11_array[c12][d358][n358];
        end
    endgenerate
    generate 
        localparam integer d359 = 23;
        for (n359 = 0; n359 < 16; n359 = n359 + 1) 
        begin: outbit359
            assign data_11[n359 + d359*16 + c12*28*16] = data_11_array[c12][d359][n359];
        end
    endgenerate
    generate 
        localparam integer d360 = 24;
        for (n360 = 0; n360 < 16; n360 = n360 + 1) 
        begin: outbit360
            assign data_11[n360 + d360*16 + c12*28*16] = data_11_array[c12][d360][n360];
        end
    endgenerate
    generate 
        localparam integer d361 = 25;
        for (n361 = 0; n361 < 16; n361 = n361 + 1) 
        begin: outbit361
            assign data_11[n361 + d361*16 + c12*28*16] = data_11_array[c12][d361][n361];
        end
    endgenerate
    generate 
        localparam integer d362 = 26;
        for (n362 = 0; n362 < 16; n362 = n362 + 1) 
        begin: outbit362
            assign data_11[n362 + d362*16 + c12*28*16] = data_11_array[c12][d362][n362];
        end
    endgenerate
    generate 
        localparam integer d363 = 27;
        for (n363 = 0; n363 < 16; n363 = n363 + 1) 
        begin: outbit363
            assign data_11[n363 + d363*16 + c12*28*16] = data_11_array[c12][d363][n363];
        end
    endgenerate
    localparam integer c13 = 13;
    generate 
        localparam integer d364 = 0;
        for (n364 = 0; n364 < 16; n364 = n364 + 1) 
        begin: outbit364
            assign data_11[n364 + d364*16 + c13*28*16] = data_11_array[c13][d364][n364];
        end
    endgenerate
    generate 
        localparam integer d365 = 1;
        for (n365 = 0; n365 < 16; n365 = n365 + 1) 
        begin: outbit365
            assign data_11[n365 + d365*16 + c13*28*16] = data_11_array[c13][d365][n365];
        end
    endgenerate
    generate 
        localparam integer d366 = 2;
        for (n366 = 0; n366 < 16; n366 = n366 + 1) 
        begin: outbit366
            assign data_11[n366 + d366*16 + c13*28*16] = data_11_array[c13][d366][n366];
        end
    endgenerate
    generate 
        localparam integer d367 = 3;
        for (n367 = 0; n367 < 16; n367 = n367 + 1) 
        begin: outbit367
            assign data_11[n367 + d367*16 + c13*28*16] = data_11_array[c13][d367][n367];
        end
    endgenerate
    generate 
        localparam integer d368 = 4;
        for (n368 = 0; n368 < 16; n368 = n368 + 1) 
        begin: outbit368
            assign data_11[n368 + d368*16 + c13*28*16] = data_11_array[c13][d368][n368];
        end
    endgenerate
    generate 
        localparam integer d369 = 5;
        for (n369 = 0; n369 < 16; n369 = n369 + 1) 
        begin: outbit369
            assign data_11[n369 + d369*16 + c13*28*16] = data_11_array[c13][d369][n369];
        end
    endgenerate
    generate 
        localparam integer d370 = 6;
        for (n370 = 0; n370 < 16; n370 = n370 + 1) 
        begin: outbit370
            assign data_11[n370 + d370*16 + c13*28*16] = data_11_array[c13][d370][n370];
        end
    endgenerate
    generate 
        localparam integer d371 = 7;
        for (n371 = 0; n371 < 16; n371 = n371 + 1) 
        begin: outbit371
            assign data_11[n371 + d371*16 + c13*28*16] = data_11_array[c13][d371][n371];
        end
    endgenerate
    generate 
        localparam integer d372 = 8;
        for (n372 = 0; n372 < 16; n372 = n372 + 1) 
        begin: outbit372
            assign data_11[n372 + d372*16 + c13*28*16] = data_11_array[c13][d372][n372];
        end
    endgenerate
    generate 
        localparam integer d373 = 9;
        for (n373 = 0; n373 < 16; n373 = n373 + 1) 
        begin: outbit373
            assign data_11[n373 + d373*16 + c13*28*16] = data_11_array[c13][d373][n373];
        end
    endgenerate
    generate 
        localparam integer d374 = 10;
        for (n374 = 0; n374 < 16; n374 = n374 + 1) 
        begin: outbit374
            assign data_11[n374 + d374*16 + c13*28*16] = data_11_array[c13][d374][n374];
        end
    endgenerate
    generate 
        localparam integer d375 = 11;
        for (n375 = 0; n375 < 16; n375 = n375 + 1) 
        begin: outbit375
            assign data_11[n375 + d375*16 + c13*28*16] = data_11_array[c13][d375][n375];
        end
    endgenerate
    generate 
        localparam integer d376 = 12;
        for (n376 = 0; n376 < 16; n376 = n376 + 1) 
        begin: outbit376
            assign data_11[n376 + d376*16 + c13*28*16] = data_11_array[c13][d376][n376];
        end
    endgenerate
    generate 
        localparam integer d377 = 13;
        for (n377 = 0; n377 < 16; n377 = n377 + 1) 
        begin: outbit377
            assign data_11[n377 + d377*16 + c13*28*16] = data_11_array[c13][d377][n377];
        end
    endgenerate
    generate 
        localparam integer d378 = 14;
        for (n378 = 0; n378 < 16; n378 = n378 + 1) 
        begin: outbit378
            assign data_11[n378 + d378*16 + c13*28*16] = data_11_array[c13][d378][n378];
        end
    endgenerate
    generate 
        localparam integer d379 = 15;
        for (n379 = 0; n379 < 16; n379 = n379 + 1) 
        begin: outbit379
            assign data_11[n379 + d379*16 + c13*28*16] = data_11_array[c13][d379][n379];
        end
    endgenerate
    generate 
        localparam integer d380 = 16;
        for (n380 = 0; n380 < 16; n380 = n380 + 1) 
        begin: outbit380
            assign data_11[n380 + d380*16 + c13*28*16] = data_11_array[c13][d380][n380];
        end
    endgenerate
    generate 
        localparam integer d381 = 17;
        for (n381 = 0; n381 < 16; n381 = n381 + 1) 
        begin: outbit381
            assign data_11[n381 + d381*16 + c13*28*16] = data_11_array[c13][d381][n381];
        end
    endgenerate
    generate 
        localparam integer d382 = 18;
        for (n382 = 0; n382 < 16; n382 = n382 + 1) 
        begin: outbit382
            assign data_11[n382 + d382*16 + c13*28*16] = data_11_array[c13][d382][n382];
        end
    endgenerate
    generate 
        localparam integer d383 = 19;
        for (n383 = 0; n383 < 16; n383 = n383 + 1) 
        begin: outbit383
            assign data_11[n383 + d383*16 + c13*28*16] = data_11_array[c13][d383][n383];
        end
    endgenerate
    generate 
        localparam integer d384 = 20;
        for (n384 = 0; n384 < 16; n384 = n384 + 1) 
        begin: outbit384
            assign data_11[n384 + d384*16 + c13*28*16] = data_11_array[c13][d384][n384];
        end
    endgenerate
    generate 
        localparam integer d385 = 21;
        for (n385 = 0; n385 < 16; n385 = n385 + 1) 
        begin: outbit385
            assign data_11[n385 + d385*16 + c13*28*16] = data_11_array[c13][d385][n385];
        end
    endgenerate
    generate 
        localparam integer d386 = 22;
        for (n386 = 0; n386 < 16; n386 = n386 + 1) 
        begin: outbit386
            assign data_11[n386 + d386*16 + c13*28*16] = data_11_array[c13][d386][n386];
        end
    endgenerate
    generate 
        localparam integer d387 = 23;
        for (n387 = 0; n387 < 16; n387 = n387 + 1) 
        begin: outbit387
            assign data_11[n387 + d387*16 + c13*28*16] = data_11_array[c13][d387][n387];
        end
    endgenerate
    generate 
        localparam integer d388 = 24;
        for (n388 = 0; n388 < 16; n388 = n388 + 1) 
        begin: outbit388
            assign data_11[n388 + d388*16 + c13*28*16] = data_11_array[c13][d388][n388];
        end
    endgenerate
    generate 
        localparam integer d389 = 25;
        for (n389 = 0; n389 < 16; n389 = n389 + 1) 
        begin: outbit389
            assign data_11[n389 + d389*16 + c13*28*16] = data_11_array[c13][d389][n389];
        end
    endgenerate
    generate 
        localparam integer d390 = 26;
        for (n390 = 0; n390 < 16; n390 = n390 + 1) 
        begin: outbit390
            assign data_11[n390 + d390*16 + c13*28*16] = data_11_array[c13][d390][n390];
        end
    endgenerate
    generate 
        localparam integer d391 = 27;
        for (n391 = 0; n391 < 16; n391 = n391 + 1) 
        begin: outbit391
            assign data_11[n391 + d391*16 + c13*28*16] = data_11_array[c13][d391][n391];
        end
    endgenerate
    localparam integer c14 = 14;
    generate 
        localparam integer d392 = 0;
        for (n392 = 0; n392 < 16; n392 = n392 + 1) 
        begin: outbit392
            assign data_11[n392 + d392*16 + c14*28*16] = data_11_array[c14][d392][n392];
        end
    endgenerate
    generate 
        localparam integer d393 = 1;
        for (n393 = 0; n393 < 16; n393 = n393 + 1) 
        begin: outbit393
            assign data_11[n393 + d393*16 + c14*28*16] = data_11_array[c14][d393][n393];
        end
    endgenerate
    generate 
        localparam integer d394 = 2;
        for (n394 = 0; n394 < 16; n394 = n394 + 1) 
        begin: outbit394
            assign data_11[n394 + d394*16 + c14*28*16] = data_11_array[c14][d394][n394];
        end
    endgenerate
    generate 
        localparam integer d395 = 3;
        for (n395 = 0; n395 < 16; n395 = n395 + 1) 
        begin: outbit395
            assign data_11[n395 + d395*16 + c14*28*16] = data_11_array[c14][d395][n395];
        end
    endgenerate
    generate 
        localparam integer d396 = 4;
        for (n396 = 0; n396 < 16; n396 = n396 + 1) 
        begin: outbit396
            assign data_11[n396 + d396*16 + c14*28*16] = data_11_array[c14][d396][n396];
        end
    endgenerate
    generate 
        localparam integer d397 = 5;
        for (n397 = 0; n397 < 16; n397 = n397 + 1) 
        begin: outbit397
            assign data_11[n397 + d397*16 + c14*28*16] = data_11_array[c14][d397][n397];
        end
    endgenerate
    generate 
        localparam integer d398 = 6;
        for (n398 = 0; n398 < 16; n398 = n398 + 1) 
        begin: outbit398
            assign data_11[n398 + d398*16 + c14*28*16] = data_11_array[c14][d398][n398];
        end
    endgenerate
    generate 
        localparam integer d399 = 7;
        for (n399 = 0; n399 < 16; n399 = n399 + 1) 
        begin: outbit399
            assign data_11[n399 + d399*16 + c14*28*16] = data_11_array[c14][d399][n399];
        end
    endgenerate
    generate 
        localparam integer d400 = 8;
        for (n400 = 0; n400 < 16; n400 = n400 + 1) 
        begin: outbit400
            assign data_11[n400 + d400*16 + c14*28*16] = data_11_array[c14][d400][n400];
        end
    endgenerate
    generate 
        localparam integer d401 = 9;
        for (n401 = 0; n401 < 16; n401 = n401 + 1) 
        begin: outbit401
            assign data_11[n401 + d401*16 + c14*28*16] = data_11_array[c14][d401][n401];
        end
    endgenerate
    generate 
        localparam integer d402 = 10;
        for (n402 = 0; n402 < 16; n402 = n402 + 1) 
        begin: outbit402
            assign data_11[n402 + d402*16 + c14*28*16] = data_11_array[c14][d402][n402];
        end
    endgenerate
    generate 
        localparam integer d403 = 11;
        for (n403 = 0; n403 < 16; n403 = n403 + 1) 
        begin: outbit403
            assign data_11[n403 + d403*16 + c14*28*16] = data_11_array[c14][d403][n403];
        end
    endgenerate
    generate 
        localparam integer d404 = 12;
        for (n404 = 0; n404 < 16; n404 = n404 + 1) 
        begin: outbit404
            assign data_11[n404 + d404*16 + c14*28*16] = data_11_array[c14][d404][n404];
        end
    endgenerate
    generate 
        localparam integer d405 = 13;
        for (n405 = 0; n405 < 16; n405 = n405 + 1) 
        begin: outbit405
            assign data_11[n405 + d405*16 + c14*28*16] = data_11_array[c14][d405][n405];
        end
    endgenerate
    generate 
        localparam integer d406 = 14;
        for (n406 = 0; n406 < 16; n406 = n406 + 1) 
        begin: outbit406
            assign data_11[n406 + d406*16 + c14*28*16] = data_11_array[c14][d406][n406];
        end
    endgenerate
    generate 
        localparam integer d407 = 15;
        for (n407 = 0; n407 < 16; n407 = n407 + 1) 
        begin: outbit407
            assign data_11[n407 + d407*16 + c14*28*16] = data_11_array[c14][d407][n407];
        end
    endgenerate
    generate 
        localparam integer d408 = 16;
        for (n408 = 0; n408 < 16; n408 = n408 + 1) 
        begin: outbit408
            assign data_11[n408 + d408*16 + c14*28*16] = data_11_array[c14][d408][n408];
        end
    endgenerate
    generate 
        localparam integer d409 = 17;
        for (n409 = 0; n409 < 16; n409 = n409 + 1) 
        begin: outbit409
            assign data_11[n409 + d409*16 + c14*28*16] = data_11_array[c14][d409][n409];
        end
    endgenerate
    generate 
        localparam integer d410 = 18;
        for (n410 = 0; n410 < 16; n410 = n410 + 1) 
        begin: outbit410
            assign data_11[n410 + d410*16 + c14*28*16] = data_11_array[c14][d410][n410];
        end
    endgenerate
    generate 
        localparam integer d411 = 19;
        for (n411 = 0; n411 < 16; n411 = n411 + 1) 
        begin: outbit411
            assign data_11[n411 + d411*16 + c14*28*16] = data_11_array[c14][d411][n411];
        end
    endgenerate
    generate 
        localparam integer d412 = 20;
        for (n412 = 0; n412 < 16; n412 = n412 + 1) 
        begin: outbit412
            assign data_11[n412 + d412*16 + c14*28*16] = data_11_array[c14][d412][n412];
        end
    endgenerate
    generate 
        localparam integer d413 = 21;
        for (n413 = 0; n413 < 16; n413 = n413 + 1) 
        begin: outbit413
            assign data_11[n413 + d413*16 + c14*28*16] = data_11_array[c14][d413][n413];
        end
    endgenerate
    generate 
        localparam integer d414 = 22;
        for (n414 = 0; n414 < 16; n414 = n414 + 1) 
        begin: outbit414
            assign data_11[n414 + d414*16 + c14*28*16] = data_11_array[c14][d414][n414];
        end
    endgenerate
    generate 
        localparam integer d415 = 23;
        for (n415 = 0; n415 < 16; n415 = n415 + 1) 
        begin: outbit415
            assign data_11[n415 + d415*16 + c14*28*16] = data_11_array[c14][d415][n415];
        end
    endgenerate
    generate 
        localparam integer d416 = 24;
        for (n416 = 0; n416 < 16; n416 = n416 + 1) 
        begin: outbit416
            assign data_11[n416 + d416*16 + c14*28*16] = data_11_array[c14][d416][n416];
        end
    endgenerate
    generate 
        localparam integer d417 = 25;
        for (n417 = 0; n417 < 16; n417 = n417 + 1) 
        begin: outbit417
            assign data_11[n417 + d417*16 + c14*28*16] = data_11_array[c14][d417][n417];
        end
    endgenerate
    generate 
        localparam integer d418 = 26;
        for (n418 = 0; n418 < 16; n418 = n418 + 1) 
        begin: outbit418
            assign data_11[n418 + d418*16 + c14*28*16] = data_11_array[c14][d418][n418];
        end
    endgenerate
    generate 
        localparam integer d419 = 27;
        for (n419 = 0; n419 < 16; n419 = n419 + 1) 
        begin: outbit419
            assign data_11[n419 + d419*16 + c14*28*16] = data_11_array[c14][d419][n419];
        end
    endgenerate
    localparam integer c15 = 15;
    generate 
        localparam integer d420 = 0;
        for (n420 = 0; n420 < 16; n420 = n420 + 1) 
        begin: outbit420
            assign data_11[n420 + d420*16 + c15*28*16] = data_11_array[c15][d420][n420];
        end
    endgenerate
    generate 
        localparam integer d421 = 1;
        for (n421 = 0; n421 < 16; n421 = n421 + 1) 
        begin: outbit421
            assign data_11[n421 + d421*16 + c15*28*16] = data_11_array[c15][d421][n421];
        end
    endgenerate
    generate 
        localparam integer d422 = 2;
        for (n422 = 0; n422 < 16; n422 = n422 + 1) 
        begin: outbit422
            assign data_11[n422 + d422*16 + c15*28*16] = data_11_array[c15][d422][n422];
        end
    endgenerate
    generate 
        localparam integer d423 = 3;
        for (n423 = 0; n423 < 16; n423 = n423 + 1) 
        begin: outbit423
            assign data_11[n423 + d423*16 + c15*28*16] = data_11_array[c15][d423][n423];
        end
    endgenerate
    generate 
        localparam integer d424 = 4;
        for (n424 = 0; n424 < 16; n424 = n424 + 1) 
        begin: outbit424
            assign data_11[n424 + d424*16 + c15*28*16] = data_11_array[c15][d424][n424];
        end
    endgenerate
    generate 
        localparam integer d425 = 5;
        for (n425 = 0; n425 < 16; n425 = n425 + 1) 
        begin: outbit425
            assign data_11[n425 + d425*16 + c15*28*16] = data_11_array[c15][d425][n425];
        end
    endgenerate
    generate 
        localparam integer d426 = 6;
        for (n426 = 0; n426 < 16; n426 = n426 + 1) 
        begin: outbit426
            assign data_11[n426 + d426*16 + c15*28*16] = data_11_array[c15][d426][n426];
        end
    endgenerate
    generate 
        localparam integer d427 = 7;
        for (n427 = 0; n427 < 16; n427 = n427 + 1) 
        begin: outbit427
            assign data_11[n427 + d427*16 + c15*28*16] = data_11_array[c15][d427][n427];
        end
    endgenerate
    generate 
        localparam integer d428 = 8;
        for (n428 = 0; n428 < 16; n428 = n428 + 1) 
        begin: outbit428
            assign data_11[n428 + d428*16 + c15*28*16] = data_11_array[c15][d428][n428];
        end
    endgenerate
    generate 
        localparam integer d429 = 9;
        for (n429 = 0; n429 < 16; n429 = n429 + 1) 
        begin: outbit429
            assign data_11[n429 + d429*16 + c15*28*16] = data_11_array[c15][d429][n429];
        end
    endgenerate
    generate 
        localparam integer d430 = 10;
        for (n430 = 0; n430 < 16; n430 = n430 + 1) 
        begin: outbit430
            assign data_11[n430 + d430*16 + c15*28*16] = data_11_array[c15][d430][n430];
        end
    endgenerate
    generate 
        localparam integer d431 = 11;
        for (n431 = 0; n431 < 16; n431 = n431 + 1) 
        begin: outbit431
            assign data_11[n431 + d431*16 + c15*28*16] = data_11_array[c15][d431][n431];
        end
    endgenerate
    generate 
        localparam integer d432 = 12;
        for (n432 = 0; n432 < 16; n432 = n432 + 1) 
        begin: outbit432
            assign data_11[n432 + d432*16 + c15*28*16] = data_11_array[c15][d432][n432];
        end
    endgenerate
    generate 
        localparam integer d433 = 13;
        for (n433 = 0; n433 < 16; n433 = n433 + 1) 
        begin: outbit433
            assign data_11[n433 + d433*16 + c15*28*16] = data_11_array[c15][d433][n433];
        end
    endgenerate
    generate 
        localparam integer d434 = 14;
        for (n434 = 0; n434 < 16; n434 = n434 + 1) 
        begin: outbit434
            assign data_11[n434 + d434*16 + c15*28*16] = data_11_array[c15][d434][n434];
        end
    endgenerate
    generate 
        localparam integer d435 = 15;
        for (n435 = 0; n435 < 16; n435 = n435 + 1) 
        begin: outbit435
            assign data_11[n435 + d435*16 + c15*28*16] = data_11_array[c15][d435][n435];
        end
    endgenerate
    generate 
        localparam integer d436 = 16;
        for (n436 = 0; n436 < 16; n436 = n436 + 1) 
        begin: outbit436
            assign data_11[n436 + d436*16 + c15*28*16] = data_11_array[c15][d436][n436];
        end
    endgenerate
    generate 
        localparam integer d437 = 17;
        for (n437 = 0; n437 < 16; n437 = n437 + 1) 
        begin: outbit437
            assign data_11[n437 + d437*16 + c15*28*16] = data_11_array[c15][d437][n437];
        end
    endgenerate
    generate 
        localparam integer d438 = 18;
        for (n438 = 0; n438 < 16; n438 = n438 + 1) 
        begin: outbit438
            assign data_11[n438 + d438*16 + c15*28*16] = data_11_array[c15][d438][n438];
        end
    endgenerate
    generate 
        localparam integer d439 = 19;
        for (n439 = 0; n439 < 16; n439 = n439 + 1) 
        begin: outbit439
            assign data_11[n439 + d439*16 + c15*28*16] = data_11_array[c15][d439][n439];
        end
    endgenerate
    generate 
        localparam integer d440 = 20;
        for (n440 = 0; n440 < 16; n440 = n440 + 1) 
        begin: outbit440
            assign data_11[n440 + d440*16 + c15*28*16] = data_11_array[c15][d440][n440];
        end
    endgenerate
    generate 
        localparam integer d441 = 21;
        for (n441 = 0; n441 < 16; n441 = n441 + 1) 
        begin: outbit441
            assign data_11[n441 + d441*16 + c15*28*16] = data_11_array[c15][d441][n441];
        end
    endgenerate
    generate 
        localparam integer d442 = 22;
        for (n442 = 0; n442 < 16; n442 = n442 + 1) 
        begin: outbit442
            assign data_11[n442 + d442*16 + c15*28*16] = data_11_array[c15][d442][n442];
        end
    endgenerate
    generate 
        localparam integer d443 = 23;
        for (n443 = 0; n443 < 16; n443 = n443 + 1) 
        begin: outbit443
            assign data_11[n443 + d443*16 + c15*28*16] = data_11_array[c15][d443][n443];
        end
    endgenerate
    generate 
        localparam integer d444 = 24;
        for (n444 = 0; n444 < 16; n444 = n444 + 1) 
        begin: outbit444
            assign data_11[n444 + d444*16 + c15*28*16] = data_11_array[c15][d444][n444];
        end
    endgenerate
    generate 
        localparam integer d445 = 25;
        for (n445 = 0; n445 < 16; n445 = n445 + 1) 
        begin: outbit445
            assign data_11[n445 + d445*16 + c15*28*16] = data_11_array[c15][d445][n445];
        end
    endgenerate
    generate 
        localparam integer d446 = 26;
        for (n446 = 0; n446 < 16; n446 = n446 + 1) 
        begin: outbit446
            assign data_11[n446 + d446*16 + c15*28*16] = data_11_array[c15][d446][n446];
        end
    endgenerate
    generate 
        localparam integer d447 = 27;
        for (n447 = 0; n447 < 16; n447 = n447 + 1) 
        begin: outbit447
            assign data_11[n447 + d447*16 + c15*28*16] = data_11_array[c15][d447][n447];
        end
    endgenerate
    localparam integer c16 = 16;
    generate 
        localparam integer d448 = 0;
        for (n448 = 0; n448 < 16; n448 = n448 + 1) 
        begin: outbit448
            assign data_11[n448 + d448*16 + c16*28*16] = data_11_array[c16][d448][n448];
        end
    endgenerate
    generate 
        localparam integer d449 = 1;
        for (n449 = 0; n449 < 16; n449 = n449 + 1) 
        begin: outbit449
            assign data_11[n449 + d449*16 + c16*28*16] = data_11_array[c16][d449][n449];
        end
    endgenerate
    generate 
        localparam integer d450 = 2;
        for (n450 = 0; n450 < 16; n450 = n450 + 1) 
        begin: outbit450
            assign data_11[n450 + d450*16 + c16*28*16] = data_11_array[c16][d450][n450];
        end
    endgenerate
    generate 
        localparam integer d451 = 3;
        for (n451 = 0; n451 < 16; n451 = n451 + 1) 
        begin: outbit451
            assign data_11[n451 + d451*16 + c16*28*16] = data_11_array[c16][d451][n451];
        end
    endgenerate
    generate 
        localparam integer d452 = 4;
        for (n452 = 0; n452 < 16; n452 = n452 + 1) 
        begin: outbit452
            assign data_11[n452 + d452*16 + c16*28*16] = data_11_array[c16][d452][n452];
        end
    endgenerate
    generate 
        localparam integer d453 = 5;
        for (n453 = 0; n453 < 16; n453 = n453 + 1) 
        begin: outbit453
            assign data_11[n453 + d453*16 + c16*28*16] = data_11_array[c16][d453][n453];
        end
    endgenerate
    generate 
        localparam integer d454 = 6;
        for (n454 = 0; n454 < 16; n454 = n454 + 1) 
        begin: outbit454
            assign data_11[n454 + d454*16 + c16*28*16] = data_11_array[c16][d454][n454];
        end
    endgenerate
    generate 
        localparam integer d455 = 7;
        for (n455 = 0; n455 < 16; n455 = n455 + 1) 
        begin: outbit455
            assign data_11[n455 + d455*16 + c16*28*16] = data_11_array[c16][d455][n455];
        end
    endgenerate
    generate 
        localparam integer d456 = 8;
        for (n456 = 0; n456 < 16; n456 = n456 + 1) 
        begin: outbit456
            assign data_11[n456 + d456*16 + c16*28*16] = data_11_array[c16][d456][n456];
        end
    endgenerate
    generate 
        localparam integer d457 = 9;
        for (n457 = 0; n457 < 16; n457 = n457 + 1) 
        begin: outbit457
            assign data_11[n457 + d457*16 + c16*28*16] = data_11_array[c16][d457][n457];
        end
    endgenerate
    generate 
        localparam integer d458 = 10;
        for (n458 = 0; n458 < 16; n458 = n458 + 1) 
        begin: outbit458
            assign data_11[n458 + d458*16 + c16*28*16] = data_11_array[c16][d458][n458];
        end
    endgenerate
    generate 
        localparam integer d459 = 11;
        for (n459 = 0; n459 < 16; n459 = n459 + 1) 
        begin: outbit459
            assign data_11[n459 + d459*16 + c16*28*16] = data_11_array[c16][d459][n459];
        end
    endgenerate
    generate 
        localparam integer d460 = 12;
        for (n460 = 0; n460 < 16; n460 = n460 + 1) 
        begin: outbit460
            assign data_11[n460 + d460*16 + c16*28*16] = data_11_array[c16][d460][n460];
        end
    endgenerate
    generate 
        localparam integer d461 = 13;
        for (n461 = 0; n461 < 16; n461 = n461 + 1) 
        begin: outbit461
            assign data_11[n461 + d461*16 + c16*28*16] = data_11_array[c16][d461][n461];
        end
    endgenerate
    generate 
        localparam integer d462 = 14;
        for (n462 = 0; n462 < 16; n462 = n462 + 1) 
        begin: outbit462
            assign data_11[n462 + d462*16 + c16*28*16] = data_11_array[c16][d462][n462];
        end
    endgenerate
    generate 
        localparam integer d463 = 15;
        for (n463 = 0; n463 < 16; n463 = n463 + 1) 
        begin: outbit463
            assign data_11[n463 + d463*16 + c16*28*16] = data_11_array[c16][d463][n463];
        end
    endgenerate
    generate 
        localparam integer d464 = 16;
        for (n464 = 0; n464 < 16; n464 = n464 + 1) 
        begin: outbit464
            assign data_11[n464 + d464*16 + c16*28*16] = data_11_array[c16][d464][n464];
        end
    endgenerate
    generate 
        localparam integer d465 = 17;
        for (n465 = 0; n465 < 16; n465 = n465 + 1) 
        begin: outbit465
            assign data_11[n465 + d465*16 + c16*28*16] = data_11_array[c16][d465][n465];
        end
    endgenerate
    generate 
        localparam integer d466 = 18;
        for (n466 = 0; n466 < 16; n466 = n466 + 1) 
        begin: outbit466
            assign data_11[n466 + d466*16 + c16*28*16] = data_11_array[c16][d466][n466];
        end
    endgenerate
    generate 
        localparam integer d467 = 19;
        for (n467 = 0; n467 < 16; n467 = n467 + 1) 
        begin: outbit467
            assign data_11[n467 + d467*16 + c16*28*16] = data_11_array[c16][d467][n467];
        end
    endgenerate
    generate 
        localparam integer d468 = 20;
        for (n468 = 0; n468 < 16; n468 = n468 + 1) 
        begin: outbit468
            assign data_11[n468 + d468*16 + c16*28*16] = data_11_array[c16][d468][n468];
        end
    endgenerate
    generate 
        localparam integer d469 = 21;
        for (n469 = 0; n469 < 16; n469 = n469 + 1) 
        begin: outbit469
            assign data_11[n469 + d469*16 + c16*28*16] = data_11_array[c16][d469][n469];
        end
    endgenerate
    generate 
        localparam integer d470 = 22;
        for (n470 = 0; n470 < 16; n470 = n470 + 1) 
        begin: outbit470
            assign data_11[n470 + d470*16 + c16*28*16] = data_11_array[c16][d470][n470];
        end
    endgenerate
    generate 
        localparam integer d471 = 23;
        for (n471 = 0; n471 < 16; n471 = n471 + 1) 
        begin: outbit471
            assign data_11[n471 + d471*16 + c16*28*16] = data_11_array[c16][d471][n471];
        end
    endgenerate
    generate 
        localparam integer d472 = 24;
        for (n472 = 0; n472 < 16; n472 = n472 + 1) 
        begin: outbit472
            assign data_11[n472 + d472*16 + c16*28*16] = data_11_array[c16][d472][n472];
        end
    endgenerate
    generate 
        localparam integer d473 = 25;
        for (n473 = 0; n473 < 16; n473 = n473 + 1) 
        begin: outbit473
            assign data_11[n473 + d473*16 + c16*28*16] = data_11_array[c16][d473][n473];
        end
    endgenerate
    generate 
        localparam integer d474 = 26;
        for (n474 = 0; n474 < 16; n474 = n474 + 1) 
        begin: outbit474
            assign data_11[n474 + d474*16 + c16*28*16] = data_11_array[c16][d474][n474];
        end
    endgenerate
    generate 
        localparam integer d475 = 27;
        for (n475 = 0; n475 < 16; n475 = n475 + 1) 
        begin: outbit475
            assign data_11[n475 + d475*16 + c16*28*16] = data_11_array[c16][d475][n475];
        end
    endgenerate
    localparam integer c17 = 17;
    generate 
        localparam integer d476 = 0;
        for (n476 = 0; n476 < 16; n476 = n476 + 1) 
        begin: outbit476
            assign data_11[n476 + d476*16 + c17*28*16] = data_11_array[c17][d476][n476];
        end
    endgenerate
    generate 
        localparam integer d477 = 1;
        for (n477 = 0; n477 < 16; n477 = n477 + 1) 
        begin: outbit477
            assign data_11[n477 + d477*16 + c17*28*16] = data_11_array[c17][d477][n477];
        end
    endgenerate
    generate 
        localparam integer d478 = 2;
        for (n478 = 0; n478 < 16; n478 = n478 + 1) 
        begin: outbit478
            assign data_11[n478 + d478*16 + c17*28*16] = data_11_array[c17][d478][n478];
        end
    endgenerate
    generate 
        localparam integer d479 = 3;
        for (n479 = 0; n479 < 16; n479 = n479 + 1) 
        begin: outbit479
            assign data_11[n479 + d479*16 + c17*28*16] = data_11_array[c17][d479][n479];
        end
    endgenerate
    generate 
        localparam integer d480 = 4;
        for (n480 = 0; n480 < 16; n480 = n480 + 1) 
        begin: outbit480
            assign data_11[n480 + d480*16 + c17*28*16] = data_11_array[c17][d480][n480];
        end
    endgenerate
    generate 
        localparam integer d481 = 5;
        for (n481 = 0; n481 < 16; n481 = n481 + 1) 
        begin: outbit481
            assign data_11[n481 + d481*16 + c17*28*16] = data_11_array[c17][d481][n481];
        end
    endgenerate
    generate 
        localparam integer d482 = 6;
        for (n482 = 0; n482 < 16; n482 = n482 + 1) 
        begin: outbit482
            assign data_11[n482 + d482*16 + c17*28*16] = data_11_array[c17][d482][n482];
        end
    endgenerate
    generate 
        localparam integer d483 = 7;
        for (n483 = 0; n483 < 16; n483 = n483 + 1) 
        begin: outbit483
            assign data_11[n483 + d483*16 + c17*28*16] = data_11_array[c17][d483][n483];
        end
    endgenerate
    generate 
        localparam integer d484 = 8;
        for (n484 = 0; n484 < 16; n484 = n484 + 1) 
        begin: outbit484
            assign data_11[n484 + d484*16 + c17*28*16] = data_11_array[c17][d484][n484];
        end
    endgenerate
    generate 
        localparam integer d485 = 9;
        for (n485 = 0; n485 < 16; n485 = n485 + 1) 
        begin: outbit485
            assign data_11[n485 + d485*16 + c17*28*16] = data_11_array[c17][d485][n485];
        end
    endgenerate
    generate 
        localparam integer d486 = 10;
        for (n486 = 0; n486 < 16; n486 = n486 + 1) 
        begin: outbit486
            assign data_11[n486 + d486*16 + c17*28*16] = data_11_array[c17][d486][n486];
        end
    endgenerate
    generate 
        localparam integer d487 = 11;
        for (n487 = 0; n487 < 16; n487 = n487 + 1) 
        begin: outbit487
            assign data_11[n487 + d487*16 + c17*28*16] = data_11_array[c17][d487][n487];
        end
    endgenerate
    generate 
        localparam integer d488 = 12;
        for (n488 = 0; n488 < 16; n488 = n488 + 1) 
        begin: outbit488
            assign data_11[n488 + d488*16 + c17*28*16] = data_11_array[c17][d488][n488];
        end
    endgenerate
    generate 
        localparam integer d489 = 13;
        for (n489 = 0; n489 < 16; n489 = n489 + 1) 
        begin: outbit489
            assign data_11[n489 + d489*16 + c17*28*16] = data_11_array[c17][d489][n489];
        end
    endgenerate
    generate 
        localparam integer d490 = 14;
        for (n490 = 0; n490 < 16; n490 = n490 + 1) 
        begin: outbit490
            assign data_11[n490 + d490*16 + c17*28*16] = data_11_array[c17][d490][n490];
        end
    endgenerate
    generate 
        localparam integer d491 = 15;
        for (n491 = 0; n491 < 16; n491 = n491 + 1) 
        begin: outbit491
            assign data_11[n491 + d491*16 + c17*28*16] = data_11_array[c17][d491][n491];
        end
    endgenerate
    generate 
        localparam integer d492 = 16;
        for (n492 = 0; n492 < 16; n492 = n492 + 1) 
        begin: outbit492
            assign data_11[n492 + d492*16 + c17*28*16] = data_11_array[c17][d492][n492];
        end
    endgenerate
    generate 
        localparam integer d493 = 17;
        for (n493 = 0; n493 < 16; n493 = n493 + 1) 
        begin: outbit493
            assign data_11[n493 + d493*16 + c17*28*16] = data_11_array[c17][d493][n493];
        end
    endgenerate
    generate 
        localparam integer d494 = 18;
        for (n494 = 0; n494 < 16; n494 = n494 + 1) 
        begin: outbit494
            assign data_11[n494 + d494*16 + c17*28*16] = data_11_array[c17][d494][n494];
        end
    endgenerate
    generate 
        localparam integer d495 = 19;
        for (n495 = 0; n495 < 16; n495 = n495 + 1) 
        begin: outbit495
            assign data_11[n495 + d495*16 + c17*28*16] = data_11_array[c17][d495][n495];
        end
    endgenerate
    generate 
        localparam integer d496 = 20;
        for (n496 = 0; n496 < 16; n496 = n496 + 1) 
        begin: outbit496
            assign data_11[n496 + d496*16 + c17*28*16] = data_11_array[c17][d496][n496];
        end
    endgenerate
    generate 
        localparam integer d497 = 21;
        for (n497 = 0; n497 < 16; n497 = n497 + 1) 
        begin: outbit497
            assign data_11[n497 + d497*16 + c17*28*16] = data_11_array[c17][d497][n497];
        end
    endgenerate
    generate 
        localparam integer d498 = 22;
        for (n498 = 0; n498 < 16; n498 = n498 + 1) 
        begin: outbit498
            assign data_11[n498 + d498*16 + c17*28*16] = data_11_array[c17][d498][n498];
        end
    endgenerate
    generate 
        localparam integer d499 = 23;
        for (n499 = 0; n499 < 16; n499 = n499 + 1) 
        begin: outbit499
            assign data_11[n499 + d499*16 + c17*28*16] = data_11_array[c17][d499][n499];
        end
    endgenerate
    generate 
        localparam integer d500 = 24;
        for (n500 = 0; n500 < 16; n500 = n500 + 1) 
        begin: outbit500
            assign data_11[n500 + d500*16 + c17*28*16] = data_11_array[c17][d500][n500];
        end
    endgenerate
    generate 
        localparam integer d501 = 25;
        for (n501 = 0; n501 < 16; n501 = n501 + 1) 
        begin: outbit501
            assign data_11[n501 + d501*16 + c17*28*16] = data_11_array[c17][d501][n501];
        end
    endgenerate
    generate 
        localparam integer d502 = 26;
        for (n502 = 0; n502 < 16; n502 = n502 + 1) 
        begin: outbit502
            assign data_11[n502 + d502*16 + c17*28*16] = data_11_array[c17][d502][n502];
        end
    endgenerate
    generate 
        localparam integer d503 = 27;
        for (n503 = 0; n503 < 16; n503 = n503 + 1) 
        begin: outbit503
            assign data_11[n503 + d503*16 + c17*28*16] = data_11_array[c17][d503][n503];
        end
    endgenerate
    localparam integer c18 = 18;
    generate 
        localparam integer d504 = 0;
        for (n504 = 0; n504 < 16; n504 = n504 + 1) 
        begin: outbit504
            assign data_11[n504 + d504*16 + c18*28*16] = data_11_array[c18][d504][n504];
        end
    endgenerate
    generate 
        localparam integer d505 = 1;
        for (n505 = 0; n505 < 16; n505 = n505 + 1) 
        begin: outbit505
            assign data_11[n505 + d505*16 + c18*28*16] = data_11_array[c18][d505][n505];
        end
    endgenerate
    generate 
        localparam integer d506 = 2;
        for (n506 = 0; n506 < 16; n506 = n506 + 1) 
        begin: outbit506
            assign data_11[n506 + d506*16 + c18*28*16] = data_11_array[c18][d506][n506];
        end
    endgenerate
    generate 
        localparam integer d507 = 3;
        for (n507 = 0; n507 < 16; n507 = n507 + 1) 
        begin: outbit507
            assign data_11[n507 + d507*16 + c18*28*16] = data_11_array[c18][d507][n507];
        end
    endgenerate
    generate 
        localparam integer d508 = 4;
        for (n508 = 0; n508 < 16; n508 = n508 + 1) 
        begin: outbit508
            assign data_11[n508 + d508*16 + c18*28*16] = data_11_array[c18][d508][n508];
        end
    endgenerate
    generate 
        localparam integer d509 = 5;
        for (n509 = 0; n509 < 16; n509 = n509 + 1) 
        begin: outbit509
            assign data_11[n509 + d509*16 + c18*28*16] = data_11_array[c18][d509][n509];
        end
    endgenerate
    generate 
        localparam integer d510 = 6;
        for (n510 = 0; n510 < 16; n510 = n510 + 1) 
        begin: outbit510
            assign data_11[n510 + d510*16 + c18*28*16] = data_11_array[c18][d510][n510];
        end
    endgenerate
    generate 
        localparam integer d511 = 7;
        for (n511 = 0; n511 < 16; n511 = n511 + 1) 
        begin: outbit511
            assign data_11[n511 + d511*16 + c18*28*16] = data_11_array[c18][d511][n511];
        end
    endgenerate
    generate 
        localparam integer d512 = 8;
        for (n512 = 0; n512 < 16; n512 = n512 + 1) 
        begin: outbit512
            assign data_11[n512 + d512*16 + c18*28*16] = data_11_array[c18][d512][n512];
        end
    endgenerate
    generate 
        localparam integer d513 = 9;
        for (n513 = 0; n513 < 16; n513 = n513 + 1) 
        begin: outbit513
            assign data_11[n513 + d513*16 + c18*28*16] = data_11_array[c18][d513][n513];
        end
    endgenerate
    generate 
        localparam integer d514 = 10;
        for (n514 = 0; n514 < 16; n514 = n514 + 1) 
        begin: outbit514
            assign data_11[n514 + d514*16 + c18*28*16] = data_11_array[c18][d514][n514];
        end
    endgenerate
    generate 
        localparam integer d515 = 11;
        for (n515 = 0; n515 < 16; n515 = n515 + 1) 
        begin: outbit515
            assign data_11[n515 + d515*16 + c18*28*16] = data_11_array[c18][d515][n515];
        end
    endgenerate
    generate 
        localparam integer d516 = 12;
        for (n516 = 0; n516 < 16; n516 = n516 + 1) 
        begin: outbit516
            assign data_11[n516 + d516*16 + c18*28*16] = data_11_array[c18][d516][n516];
        end
    endgenerate
    generate 
        localparam integer d517 = 13;
        for (n517 = 0; n517 < 16; n517 = n517 + 1) 
        begin: outbit517
            assign data_11[n517 + d517*16 + c18*28*16] = data_11_array[c18][d517][n517];
        end
    endgenerate
    generate 
        localparam integer d518 = 14;
        for (n518 = 0; n518 < 16; n518 = n518 + 1) 
        begin: outbit518
            assign data_11[n518 + d518*16 + c18*28*16] = data_11_array[c18][d518][n518];
        end
    endgenerate
    generate 
        localparam integer d519 = 15;
        for (n519 = 0; n519 < 16; n519 = n519 + 1) 
        begin: outbit519
            assign data_11[n519 + d519*16 + c18*28*16] = data_11_array[c18][d519][n519];
        end
    endgenerate
    generate 
        localparam integer d520 = 16;
        for (n520 = 0; n520 < 16; n520 = n520 + 1) 
        begin: outbit520
            assign data_11[n520 + d520*16 + c18*28*16] = data_11_array[c18][d520][n520];
        end
    endgenerate
    generate 
        localparam integer d521 = 17;
        for (n521 = 0; n521 < 16; n521 = n521 + 1) 
        begin: outbit521
            assign data_11[n521 + d521*16 + c18*28*16] = data_11_array[c18][d521][n521];
        end
    endgenerate
    generate 
        localparam integer d522 = 18;
        for (n522 = 0; n522 < 16; n522 = n522 + 1) 
        begin: outbit522
            assign data_11[n522 + d522*16 + c18*28*16] = data_11_array[c18][d522][n522];
        end
    endgenerate
    generate 
        localparam integer d523 = 19;
        for (n523 = 0; n523 < 16; n523 = n523 + 1) 
        begin: outbit523
            assign data_11[n523 + d523*16 + c18*28*16] = data_11_array[c18][d523][n523];
        end
    endgenerate
    generate 
        localparam integer d524 = 20;
        for (n524 = 0; n524 < 16; n524 = n524 + 1) 
        begin: outbit524
            assign data_11[n524 + d524*16 + c18*28*16] = data_11_array[c18][d524][n524];
        end
    endgenerate
    generate 
        localparam integer d525 = 21;
        for (n525 = 0; n525 < 16; n525 = n525 + 1) 
        begin: outbit525
            assign data_11[n525 + d525*16 + c18*28*16] = data_11_array[c18][d525][n525];
        end
    endgenerate
    generate 
        localparam integer d526 = 22;
        for (n526 = 0; n526 < 16; n526 = n526 + 1) 
        begin: outbit526
            assign data_11[n526 + d526*16 + c18*28*16] = data_11_array[c18][d526][n526];
        end
    endgenerate
    generate 
        localparam integer d527 = 23;
        for (n527 = 0; n527 < 16; n527 = n527 + 1) 
        begin: outbit527
            assign data_11[n527 + d527*16 + c18*28*16] = data_11_array[c18][d527][n527];
        end
    endgenerate
    generate 
        localparam integer d528 = 24;
        for (n528 = 0; n528 < 16; n528 = n528 + 1) 
        begin: outbit528
            assign data_11[n528 + d528*16 + c18*28*16] = data_11_array[c18][d528][n528];
        end
    endgenerate
    generate 
        localparam integer d529 = 25;
        for (n529 = 0; n529 < 16; n529 = n529 + 1) 
        begin: outbit529
            assign data_11[n529 + d529*16 + c18*28*16] = data_11_array[c18][d529][n529];
        end
    endgenerate
    generate 
        localparam integer d530 = 26;
        for (n530 = 0; n530 < 16; n530 = n530 + 1) 
        begin: outbit530
            assign data_11[n530 + d530*16 + c18*28*16] = data_11_array[c18][d530][n530];
        end
    endgenerate
    generate 
        localparam integer d531 = 27;
        for (n531 = 0; n531 < 16; n531 = n531 + 1) 
        begin: outbit531
            assign data_11[n531 + d531*16 + c18*28*16] = data_11_array[c18][d531][n531];
        end
    endgenerate
    localparam integer c19 = 19;
    generate 
        localparam integer d532 = 0;
        for (n532 = 0; n532 < 16; n532 = n532 + 1) 
        begin: outbit532
            assign data_11[n532 + d532*16 + c19*28*16] = data_11_array[c19][d532][n532];
        end
    endgenerate
    generate 
        localparam integer d533 = 1;
        for (n533 = 0; n533 < 16; n533 = n533 + 1) 
        begin: outbit533
            assign data_11[n533 + d533*16 + c19*28*16] = data_11_array[c19][d533][n533];
        end
    endgenerate
    generate 
        localparam integer d534 = 2;
        for (n534 = 0; n534 < 16; n534 = n534 + 1) 
        begin: outbit534
            assign data_11[n534 + d534*16 + c19*28*16] = data_11_array[c19][d534][n534];
        end
    endgenerate
    generate 
        localparam integer d535 = 3;
        for (n535 = 0; n535 < 16; n535 = n535 + 1) 
        begin: outbit535
            assign data_11[n535 + d535*16 + c19*28*16] = data_11_array[c19][d535][n535];
        end
    endgenerate
    generate 
        localparam integer d536 = 4;
        for (n536 = 0; n536 < 16; n536 = n536 + 1) 
        begin: outbit536
            assign data_11[n536 + d536*16 + c19*28*16] = data_11_array[c19][d536][n536];
        end
    endgenerate
    generate 
        localparam integer d537 = 5;
        for (n537 = 0; n537 < 16; n537 = n537 + 1) 
        begin: outbit537
            assign data_11[n537 + d537*16 + c19*28*16] = data_11_array[c19][d537][n537];
        end
    endgenerate
    generate 
        localparam integer d538 = 6;
        for (n538 = 0; n538 < 16; n538 = n538 + 1) 
        begin: outbit538
            assign data_11[n538 + d538*16 + c19*28*16] = data_11_array[c19][d538][n538];
        end
    endgenerate
    generate 
        localparam integer d539 = 7;
        for (n539 = 0; n539 < 16; n539 = n539 + 1) 
        begin: outbit539
            assign data_11[n539 + d539*16 + c19*28*16] = data_11_array[c19][d539][n539];
        end
    endgenerate
    generate 
        localparam integer d540 = 8;
        for (n540 = 0; n540 < 16; n540 = n540 + 1) 
        begin: outbit540
            assign data_11[n540 + d540*16 + c19*28*16] = data_11_array[c19][d540][n540];
        end
    endgenerate
    generate 
        localparam integer d541 = 9;
        for (n541 = 0; n541 < 16; n541 = n541 + 1) 
        begin: outbit541
            assign data_11[n541 + d541*16 + c19*28*16] = data_11_array[c19][d541][n541];
        end
    endgenerate
    generate 
        localparam integer d542 = 10;
        for (n542 = 0; n542 < 16; n542 = n542 + 1) 
        begin: outbit542
            assign data_11[n542 + d542*16 + c19*28*16] = data_11_array[c19][d542][n542];
        end
    endgenerate
    generate 
        localparam integer d543 = 11;
        for (n543 = 0; n543 < 16; n543 = n543 + 1) 
        begin: outbit543
            assign data_11[n543 + d543*16 + c19*28*16] = data_11_array[c19][d543][n543];
        end
    endgenerate
    generate 
        localparam integer d544 = 12;
        for (n544 = 0; n544 < 16; n544 = n544 + 1) 
        begin: outbit544
            assign data_11[n544 + d544*16 + c19*28*16] = data_11_array[c19][d544][n544];
        end
    endgenerate
    generate 
        localparam integer d545 = 13;
        for (n545 = 0; n545 < 16; n545 = n545 + 1) 
        begin: outbit545
            assign data_11[n545 + d545*16 + c19*28*16] = data_11_array[c19][d545][n545];
        end
    endgenerate
    generate 
        localparam integer d546 = 14;
        for (n546 = 0; n546 < 16; n546 = n546 + 1) 
        begin: outbit546
            assign data_11[n546 + d546*16 + c19*28*16] = data_11_array[c19][d546][n546];
        end
    endgenerate
    generate 
        localparam integer d547 = 15;
        for (n547 = 0; n547 < 16; n547 = n547 + 1) 
        begin: outbit547
            assign data_11[n547 + d547*16 + c19*28*16] = data_11_array[c19][d547][n547];
        end
    endgenerate
    generate 
        localparam integer d548 = 16;
        for (n548 = 0; n548 < 16; n548 = n548 + 1) 
        begin: outbit548
            assign data_11[n548 + d548*16 + c19*28*16] = data_11_array[c19][d548][n548];
        end
    endgenerate
    generate 
        localparam integer d549 = 17;
        for (n549 = 0; n549 < 16; n549 = n549 + 1) 
        begin: outbit549
            assign data_11[n549 + d549*16 + c19*28*16] = data_11_array[c19][d549][n549];
        end
    endgenerate
    generate 
        localparam integer d550 = 18;
        for (n550 = 0; n550 < 16; n550 = n550 + 1) 
        begin: outbit550
            assign data_11[n550 + d550*16 + c19*28*16] = data_11_array[c19][d550][n550];
        end
    endgenerate
    generate 
        localparam integer d551 = 19;
        for (n551 = 0; n551 < 16; n551 = n551 + 1) 
        begin: outbit551
            assign data_11[n551 + d551*16 + c19*28*16] = data_11_array[c19][d551][n551];
        end
    endgenerate
    generate 
        localparam integer d552 = 20;
        for (n552 = 0; n552 < 16; n552 = n552 + 1) 
        begin: outbit552
            assign data_11[n552 + d552*16 + c19*28*16] = data_11_array[c19][d552][n552];
        end
    endgenerate
    generate 
        localparam integer d553 = 21;
        for (n553 = 0; n553 < 16; n553 = n553 + 1) 
        begin: outbit553
            assign data_11[n553 + d553*16 + c19*28*16] = data_11_array[c19][d553][n553];
        end
    endgenerate
    generate 
        localparam integer d554 = 22;
        for (n554 = 0; n554 < 16; n554 = n554 + 1) 
        begin: outbit554
            assign data_11[n554 + d554*16 + c19*28*16] = data_11_array[c19][d554][n554];
        end
    endgenerate
    generate 
        localparam integer d555 = 23;
        for (n555 = 0; n555 < 16; n555 = n555 + 1) 
        begin: outbit555
            assign data_11[n555 + d555*16 + c19*28*16] = data_11_array[c19][d555][n555];
        end
    endgenerate
    generate 
        localparam integer d556 = 24;
        for (n556 = 0; n556 < 16; n556 = n556 + 1) 
        begin: outbit556
            assign data_11[n556 + d556*16 + c19*28*16] = data_11_array[c19][d556][n556];
        end
    endgenerate
    generate 
        localparam integer d557 = 25;
        for (n557 = 0; n557 < 16; n557 = n557 + 1) 
        begin: outbit557
            assign data_11[n557 + d557*16 + c19*28*16] = data_11_array[c19][d557][n557];
        end
    endgenerate
    generate 
        localparam integer d558 = 26;
        for (n558 = 0; n558 < 16; n558 = n558 + 1) 
        begin: outbit558
            assign data_11[n558 + d558*16 + c19*28*16] = data_11_array[c19][d558][n558];
        end
    endgenerate
    generate 
        localparam integer d559 = 27;
        for (n559 = 0; n559 < 16; n559 = n559 + 1) 
        begin: outbit559
            assign data_11[n559 + d559*16 + c19*28*16] = data_11_array[c19][d559][n559];
        end
    endgenerate
    localparam integer c20 = 20;
    generate 
        localparam integer d560 = 0;
        for (n560 = 0; n560 < 16; n560 = n560 + 1) 
        begin: outbit560
            assign data_11[n560 + d560*16 + c20*28*16] = data_11_array[c20][d560][n560];
        end
    endgenerate
    generate 
        localparam integer d561 = 1;
        for (n561 = 0; n561 < 16; n561 = n561 + 1) 
        begin: outbit561
            assign data_11[n561 + d561*16 + c20*28*16] = data_11_array[c20][d561][n561];
        end
    endgenerate
    generate 
        localparam integer d562 = 2;
        for (n562 = 0; n562 < 16; n562 = n562 + 1) 
        begin: outbit562
            assign data_11[n562 + d562*16 + c20*28*16] = data_11_array[c20][d562][n562];
        end
    endgenerate
    generate 
        localparam integer d563 = 3;
        for (n563 = 0; n563 < 16; n563 = n563 + 1) 
        begin: outbit563
            assign data_11[n563 + d563*16 + c20*28*16] = data_11_array[c20][d563][n563];
        end
    endgenerate
    generate 
        localparam integer d564 = 4;
        for (n564 = 0; n564 < 16; n564 = n564 + 1) 
        begin: outbit564
            assign data_11[n564 + d564*16 + c20*28*16] = data_11_array[c20][d564][n564];
        end
    endgenerate
    generate 
        localparam integer d565 = 5;
        for (n565 = 0; n565 < 16; n565 = n565 + 1) 
        begin: outbit565
            assign data_11[n565 + d565*16 + c20*28*16] = data_11_array[c20][d565][n565];
        end
    endgenerate
    generate 
        localparam integer d566 = 6;
        for (n566 = 0; n566 < 16; n566 = n566 + 1) 
        begin: outbit566
            assign data_11[n566 + d566*16 + c20*28*16] = data_11_array[c20][d566][n566];
        end
    endgenerate
    generate 
        localparam integer d567 = 7;
        for (n567 = 0; n567 < 16; n567 = n567 + 1) 
        begin: outbit567
            assign data_11[n567 + d567*16 + c20*28*16] = data_11_array[c20][d567][n567];
        end
    endgenerate
    generate 
        localparam integer d568 = 8;
        for (n568 = 0; n568 < 16; n568 = n568 + 1) 
        begin: outbit568
            assign data_11[n568 + d568*16 + c20*28*16] = data_11_array[c20][d568][n568];
        end
    endgenerate
    generate 
        localparam integer d569 = 9;
        for (n569 = 0; n569 < 16; n569 = n569 + 1) 
        begin: outbit569
            assign data_11[n569 + d569*16 + c20*28*16] = data_11_array[c20][d569][n569];
        end
    endgenerate
    generate 
        localparam integer d570 = 10;
        for (n570 = 0; n570 < 16; n570 = n570 + 1) 
        begin: outbit570
            assign data_11[n570 + d570*16 + c20*28*16] = data_11_array[c20][d570][n570];
        end
    endgenerate
    generate 
        localparam integer d571 = 11;
        for (n571 = 0; n571 < 16; n571 = n571 + 1) 
        begin: outbit571
            assign data_11[n571 + d571*16 + c20*28*16] = data_11_array[c20][d571][n571];
        end
    endgenerate
    generate 
        localparam integer d572 = 12;
        for (n572 = 0; n572 < 16; n572 = n572 + 1) 
        begin: outbit572
            assign data_11[n572 + d572*16 + c20*28*16] = data_11_array[c20][d572][n572];
        end
    endgenerate
    generate 
        localparam integer d573 = 13;
        for (n573 = 0; n573 < 16; n573 = n573 + 1) 
        begin: outbit573
            assign data_11[n573 + d573*16 + c20*28*16] = data_11_array[c20][d573][n573];
        end
    endgenerate
    generate 
        localparam integer d574 = 14;
        for (n574 = 0; n574 < 16; n574 = n574 + 1) 
        begin: outbit574
            assign data_11[n574 + d574*16 + c20*28*16] = data_11_array[c20][d574][n574];
        end
    endgenerate
    generate 
        localparam integer d575 = 15;
        for (n575 = 0; n575 < 16; n575 = n575 + 1) 
        begin: outbit575
            assign data_11[n575 + d575*16 + c20*28*16] = data_11_array[c20][d575][n575];
        end
    endgenerate
    generate 
        localparam integer d576 = 16;
        for (n576 = 0; n576 < 16; n576 = n576 + 1) 
        begin: outbit576
            assign data_11[n576 + d576*16 + c20*28*16] = data_11_array[c20][d576][n576];
        end
    endgenerate
    generate 
        localparam integer d577 = 17;
        for (n577 = 0; n577 < 16; n577 = n577 + 1) 
        begin: outbit577
            assign data_11[n577 + d577*16 + c20*28*16] = data_11_array[c20][d577][n577];
        end
    endgenerate
    generate 
        localparam integer d578 = 18;
        for (n578 = 0; n578 < 16; n578 = n578 + 1) 
        begin: outbit578
            assign data_11[n578 + d578*16 + c20*28*16] = data_11_array[c20][d578][n578];
        end
    endgenerate
    generate 
        localparam integer d579 = 19;
        for (n579 = 0; n579 < 16; n579 = n579 + 1) 
        begin: outbit579
            assign data_11[n579 + d579*16 + c20*28*16] = data_11_array[c20][d579][n579];
        end
    endgenerate
    generate 
        localparam integer d580 = 20;
        for (n580 = 0; n580 < 16; n580 = n580 + 1) 
        begin: outbit580
            assign data_11[n580 + d580*16 + c20*28*16] = data_11_array[c20][d580][n580];
        end
    endgenerate
    generate 
        localparam integer d581 = 21;
        for (n581 = 0; n581 < 16; n581 = n581 + 1) 
        begin: outbit581
            assign data_11[n581 + d581*16 + c20*28*16] = data_11_array[c20][d581][n581];
        end
    endgenerate
    generate 
        localparam integer d582 = 22;
        for (n582 = 0; n582 < 16; n582 = n582 + 1) 
        begin: outbit582
            assign data_11[n582 + d582*16 + c20*28*16] = data_11_array[c20][d582][n582];
        end
    endgenerate
    generate 
        localparam integer d583 = 23;
        for (n583 = 0; n583 < 16; n583 = n583 + 1) 
        begin: outbit583
            assign data_11[n583 + d583*16 + c20*28*16] = data_11_array[c20][d583][n583];
        end
    endgenerate
    generate 
        localparam integer d584 = 24;
        for (n584 = 0; n584 < 16; n584 = n584 + 1) 
        begin: outbit584
            assign data_11[n584 + d584*16 + c20*28*16] = data_11_array[c20][d584][n584];
        end
    endgenerate
    generate 
        localparam integer d585 = 25;
        for (n585 = 0; n585 < 16; n585 = n585 + 1) 
        begin: outbit585
            assign data_11[n585 + d585*16 + c20*28*16] = data_11_array[c20][d585][n585];
        end
    endgenerate
    generate 
        localparam integer d586 = 26;
        for (n586 = 0; n586 < 16; n586 = n586 + 1) 
        begin: outbit586
            assign data_11[n586 + d586*16 + c20*28*16] = data_11_array[c20][d586][n586];
        end
    endgenerate
    generate 
        localparam integer d587 = 27;
        for (n587 = 0; n587 < 16; n587 = n587 + 1) 
        begin: outbit587
            assign data_11[n587 + d587*16 + c20*28*16] = data_11_array[c20][d587][n587];
        end
    endgenerate
    localparam integer c21 = 21;
    generate 
        localparam integer d588 = 0;
        for (n588 = 0; n588 < 16; n588 = n588 + 1) 
        begin: outbit588
            assign data_11[n588 + d588*16 + c21*28*16] = data_11_array[c21][d588][n588];
        end
    endgenerate
    generate 
        localparam integer d589 = 1;
        for (n589 = 0; n589 < 16; n589 = n589 + 1) 
        begin: outbit589
            assign data_11[n589 + d589*16 + c21*28*16] = data_11_array[c21][d589][n589];
        end
    endgenerate
    generate 
        localparam integer d590 = 2;
        for (n590 = 0; n590 < 16; n590 = n590 + 1) 
        begin: outbit590
            assign data_11[n590 + d590*16 + c21*28*16] = data_11_array[c21][d590][n590];
        end
    endgenerate
    generate 
        localparam integer d591 = 3;
        for (n591 = 0; n591 < 16; n591 = n591 + 1) 
        begin: outbit591
            assign data_11[n591 + d591*16 + c21*28*16] = data_11_array[c21][d591][n591];
        end
    endgenerate
    generate 
        localparam integer d592 = 4;
        for (n592 = 0; n592 < 16; n592 = n592 + 1) 
        begin: outbit592
            assign data_11[n592 + d592*16 + c21*28*16] = data_11_array[c21][d592][n592];
        end
    endgenerate
    generate 
        localparam integer d593 = 5;
        for (n593 = 0; n593 < 16; n593 = n593 + 1) 
        begin: outbit593
            assign data_11[n593 + d593*16 + c21*28*16] = data_11_array[c21][d593][n593];
        end
    endgenerate
    generate 
        localparam integer d594 = 6;
        for (n594 = 0; n594 < 16; n594 = n594 + 1) 
        begin: outbit594
            assign data_11[n594 + d594*16 + c21*28*16] = data_11_array[c21][d594][n594];
        end
    endgenerate
    generate 
        localparam integer d595 = 7;
        for (n595 = 0; n595 < 16; n595 = n595 + 1) 
        begin: outbit595
            assign data_11[n595 + d595*16 + c21*28*16] = data_11_array[c21][d595][n595];
        end
    endgenerate
    generate 
        localparam integer d596 = 8;
        for (n596 = 0; n596 < 16; n596 = n596 + 1) 
        begin: outbit596
            assign data_11[n596 + d596*16 + c21*28*16] = data_11_array[c21][d596][n596];
        end
    endgenerate
    generate 
        localparam integer d597 = 9;
        for (n597 = 0; n597 < 16; n597 = n597 + 1) 
        begin: outbit597
            assign data_11[n597 + d597*16 + c21*28*16] = data_11_array[c21][d597][n597];
        end
    endgenerate
    generate 
        localparam integer d598 = 10;
        for (n598 = 0; n598 < 16; n598 = n598 + 1) 
        begin: outbit598
            assign data_11[n598 + d598*16 + c21*28*16] = data_11_array[c21][d598][n598];
        end
    endgenerate
    generate 
        localparam integer d599 = 11;
        for (n599 = 0; n599 < 16; n599 = n599 + 1) 
        begin: outbit599
            assign data_11[n599 + d599*16 + c21*28*16] = data_11_array[c21][d599][n599];
        end
    endgenerate
    generate 
        localparam integer d600 = 12;
        for (n600 = 0; n600 < 16; n600 = n600 + 1) 
        begin: outbit600
            assign data_11[n600 + d600*16 + c21*28*16] = data_11_array[c21][d600][n600];
        end
    endgenerate
    generate 
        localparam integer d601 = 13;
        for (n601 = 0; n601 < 16; n601 = n601 + 1) 
        begin: outbit601
            assign data_11[n601 + d601*16 + c21*28*16] = data_11_array[c21][d601][n601];
        end
    endgenerate
    generate 
        localparam integer d602 = 14;
        for (n602 = 0; n602 < 16; n602 = n602 + 1) 
        begin: outbit602
            assign data_11[n602 + d602*16 + c21*28*16] = data_11_array[c21][d602][n602];
        end
    endgenerate
    generate 
        localparam integer d603 = 15;
        for (n603 = 0; n603 < 16; n603 = n603 + 1) 
        begin: outbit603
            assign data_11[n603 + d603*16 + c21*28*16] = data_11_array[c21][d603][n603];
        end
    endgenerate
    generate 
        localparam integer d604 = 16;
        for (n604 = 0; n604 < 16; n604 = n604 + 1) 
        begin: outbit604
            assign data_11[n604 + d604*16 + c21*28*16] = data_11_array[c21][d604][n604];
        end
    endgenerate
    generate 
        localparam integer d605 = 17;
        for (n605 = 0; n605 < 16; n605 = n605 + 1) 
        begin: outbit605
            assign data_11[n605 + d605*16 + c21*28*16] = data_11_array[c21][d605][n605];
        end
    endgenerate
    generate 
        localparam integer d606 = 18;
        for (n606 = 0; n606 < 16; n606 = n606 + 1) 
        begin: outbit606
            assign data_11[n606 + d606*16 + c21*28*16] = data_11_array[c21][d606][n606];
        end
    endgenerate
    generate 
        localparam integer d607 = 19;
        for (n607 = 0; n607 < 16; n607 = n607 + 1) 
        begin: outbit607
            assign data_11[n607 + d607*16 + c21*28*16] = data_11_array[c21][d607][n607];
        end
    endgenerate
    generate 
        localparam integer d608 = 20;
        for (n608 = 0; n608 < 16; n608 = n608 + 1) 
        begin: outbit608
            assign data_11[n608 + d608*16 + c21*28*16] = data_11_array[c21][d608][n608];
        end
    endgenerate
    generate 
        localparam integer d609 = 21;
        for (n609 = 0; n609 < 16; n609 = n609 + 1) 
        begin: outbit609
            assign data_11[n609 + d609*16 + c21*28*16] = data_11_array[c21][d609][n609];
        end
    endgenerate
    generate 
        localparam integer d610 = 22;
        for (n610 = 0; n610 < 16; n610 = n610 + 1) 
        begin: outbit610
            assign data_11[n610 + d610*16 + c21*28*16] = data_11_array[c21][d610][n610];
        end
    endgenerate
    generate 
        localparam integer d611 = 23;
        for (n611 = 0; n611 < 16; n611 = n611 + 1) 
        begin: outbit611
            assign data_11[n611 + d611*16 + c21*28*16] = data_11_array[c21][d611][n611];
        end
    endgenerate
    generate 
        localparam integer d612 = 24;
        for (n612 = 0; n612 < 16; n612 = n612 + 1) 
        begin: outbit612
            assign data_11[n612 + d612*16 + c21*28*16] = data_11_array[c21][d612][n612];
        end
    endgenerate
    generate 
        localparam integer d613 = 25;
        for (n613 = 0; n613 < 16; n613 = n613 + 1) 
        begin: outbit613
            assign data_11[n613 + d613*16 + c21*28*16] = data_11_array[c21][d613][n613];
        end
    endgenerate
    generate 
        localparam integer d614 = 26;
        for (n614 = 0; n614 < 16; n614 = n614 + 1) 
        begin: outbit614
            assign data_11[n614 + d614*16 + c21*28*16] = data_11_array[c21][d614][n614];
        end
    endgenerate
    generate 
        localparam integer d615 = 27;
        for (n615 = 0; n615 < 16; n615 = n615 + 1) 
        begin: outbit615
            assign data_11[n615 + d615*16 + c21*28*16] = data_11_array[c21][d615][n615];
        end
    endgenerate
    localparam integer c22 = 22;
    generate 
        localparam integer d616 = 0;
        for (n616 = 0; n616 < 16; n616 = n616 + 1) 
        begin: outbit616
            assign data_11[n616 + d616*16 + c22*28*16] = data_11_array[c22][d616][n616];
        end
    endgenerate
    generate 
        localparam integer d617 = 1;
        for (n617 = 0; n617 < 16; n617 = n617 + 1) 
        begin: outbit617
            assign data_11[n617 + d617*16 + c22*28*16] = data_11_array[c22][d617][n617];
        end
    endgenerate
    generate 
        localparam integer d618 = 2;
        for (n618 = 0; n618 < 16; n618 = n618 + 1) 
        begin: outbit618
            assign data_11[n618 + d618*16 + c22*28*16] = data_11_array[c22][d618][n618];
        end
    endgenerate
    generate 
        localparam integer d619 = 3;
        for (n619 = 0; n619 < 16; n619 = n619 + 1) 
        begin: outbit619
            assign data_11[n619 + d619*16 + c22*28*16] = data_11_array[c22][d619][n619];
        end
    endgenerate
    generate 
        localparam integer d620 = 4;
        for (n620 = 0; n620 < 16; n620 = n620 + 1) 
        begin: outbit620
            assign data_11[n620 + d620*16 + c22*28*16] = data_11_array[c22][d620][n620];
        end
    endgenerate
    generate 
        localparam integer d621 = 5;
        for (n621 = 0; n621 < 16; n621 = n621 + 1) 
        begin: outbit621
            assign data_11[n621 + d621*16 + c22*28*16] = data_11_array[c22][d621][n621];
        end
    endgenerate
    generate 
        localparam integer d622 = 6;
        for (n622 = 0; n622 < 16; n622 = n622 + 1) 
        begin: outbit622
            assign data_11[n622 + d622*16 + c22*28*16] = data_11_array[c22][d622][n622];
        end
    endgenerate
    generate 
        localparam integer d623 = 7;
        for (n623 = 0; n623 < 16; n623 = n623 + 1) 
        begin: outbit623
            assign data_11[n623 + d623*16 + c22*28*16] = data_11_array[c22][d623][n623];
        end
    endgenerate
    generate 
        localparam integer d624 = 8;
        for (n624 = 0; n624 < 16; n624 = n624 + 1) 
        begin: outbit624
            assign data_11[n624 + d624*16 + c22*28*16] = data_11_array[c22][d624][n624];
        end
    endgenerate
    generate 
        localparam integer d625 = 9;
        for (n625 = 0; n625 < 16; n625 = n625 + 1) 
        begin: outbit625
            assign data_11[n625 + d625*16 + c22*28*16] = data_11_array[c22][d625][n625];
        end
    endgenerate
    generate 
        localparam integer d626 = 10;
        for (n626 = 0; n626 < 16; n626 = n626 + 1) 
        begin: outbit626
            assign data_11[n626 + d626*16 + c22*28*16] = data_11_array[c22][d626][n626];
        end
    endgenerate
    generate 
        localparam integer d627 = 11;
        for (n627 = 0; n627 < 16; n627 = n627 + 1) 
        begin: outbit627
            assign data_11[n627 + d627*16 + c22*28*16] = data_11_array[c22][d627][n627];
        end
    endgenerate
    generate 
        localparam integer d628 = 12;
        for (n628 = 0; n628 < 16; n628 = n628 + 1) 
        begin: outbit628
            assign data_11[n628 + d628*16 + c22*28*16] = data_11_array[c22][d628][n628];
        end
    endgenerate
    generate 
        localparam integer d629 = 13;
        for (n629 = 0; n629 < 16; n629 = n629 + 1) 
        begin: outbit629
            assign data_11[n629 + d629*16 + c22*28*16] = data_11_array[c22][d629][n629];
        end
    endgenerate
    generate 
        localparam integer d630 = 14;
        for (n630 = 0; n630 < 16; n630 = n630 + 1) 
        begin: outbit630
            assign data_11[n630 + d630*16 + c22*28*16] = data_11_array[c22][d630][n630];
        end
    endgenerate
    generate 
        localparam integer d631 = 15;
        for (n631 = 0; n631 < 16; n631 = n631 + 1) 
        begin: outbit631
            assign data_11[n631 + d631*16 + c22*28*16] = data_11_array[c22][d631][n631];
        end
    endgenerate
    generate 
        localparam integer d632 = 16;
        for (n632 = 0; n632 < 16; n632 = n632 + 1) 
        begin: outbit632
            assign data_11[n632 + d632*16 + c22*28*16] = data_11_array[c22][d632][n632];
        end
    endgenerate
    generate 
        localparam integer d633 = 17;
        for (n633 = 0; n633 < 16; n633 = n633 + 1) 
        begin: outbit633
            assign data_11[n633 + d633*16 + c22*28*16] = data_11_array[c22][d633][n633];
        end
    endgenerate
    generate 
        localparam integer d634 = 18;
        for (n634 = 0; n634 < 16; n634 = n634 + 1) 
        begin: outbit634
            assign data_11[n634 + d634*16 + c22*28*16] = data_11_array[c22][d634][n634];
        end
    endgenerate
    generate 
        localparam integer d635 = 19;
        for (n635 = 0; n635 < 16; n635 = n635 + 1) 
        begin: outbit635
            assign data_11[n635 + d635*16 + c22*28*16] = data_11_array[c22][d635][n635];
        end
    endgenerate
    generate 
        localparam integer d636 = 20;
        for (n636 = 0; n636 < 16; n636 = n636 + 1) 
        begin: outbit636
            assign data_11[n636 + d636*16 + c22*28*16] = data_11_array[c22][d636][n636];
        end
    endgenerate
    generate 
        localparam integer d637 = 21;
        for (n637 = 0; n637 < 16; n637 = n637 + 1) 
        begin: outbit637
            assign data_11[n637 + d637*16 + c22*28*16] = data_11_array[c22][d637][n637];
        end
    endgenerate
    generate 
        localparam integer d638 = 22;
        for (n638 = 0; n638 < 16; n638 = n638 + 1) 
        begin: outbit638
            assign data_11[n638 + d638*16 + c22*28*16] = data_11_array[c22][d638][n638];
        end
    endgenerate
    generate 
        localparam integer d639 = 23;
        for (n639 = 0; n639 < 16; n639 = n639 + 1) 
        begin: outbit639
            assign data_11[n639 + d639*16 + c22*28*16] = data_11_array[c22][d639][n639];
        end
    endgenerate
    generate 
        localparam integer d640 = 24;
        for (n640 = 0; n640 < 16; n640 = n640 + 1) 
        begin: outbit640
            assign data_11[n640 + d640*16 + c22*28*16] = data_11_array[c22][d640][n640];
        end
    endgenerate
    generate 
        localparam integer d641 = 25;
        for (n641 = 0; n641 < 16; n641 = n641 + 1) 
        begin: outbit641
            assign data_11[n641 + d641*16 + c22*28*16] = data_11_array[c22][d641][n641];
        end
    endgenerate
    generate 
        localparam integer d642 = 26;
        for (n642 = 0; n642 < 16; n642 = n642 + 1) 
        begin: outbit642
            assign data_11[n642 + d642*16 + c22*28*16] = data_11_array[c22][d642][n642];
        end
    endgenerate
    generate 
        localparam integer d643 = 27;
        for (n643 = 0; n643 < 16; n643 = n643 + 1) 
        begin: outbit643
            assign data_11[n643 + d643*16 + c22*28*16] = data_11_array[c22][d643][n643];
        end
    endgenerate
    localparam integer c23 = 23;
    generate 
        localparam integer d644 = 0;
        for (n644 = 0; n644 < 16; n644 = n644 + 1) 
        begin: outbit644
            assign data_11[n644 + d644*16 + c23*28*16] = data_11_array[c23][d644][n644];
        end
    endgenerate
    generate 
        localparam integer d645 = 1;
        for (n645 = 0; n645 < 16; n645 = n645 + 1) 
        begin: outbit645
            assign data_11[n645 + d645*16 + c23*28*16] = data_11_array[c23][d645][n645];
        end
    endgenerate
    generate 
        localparam integer d646 = 2;
        for (n646 = 0; n646 < 16; n646 = n646 + 1) 
        begin: outbit646
            assign data_11[n646 + d646*16 + c23*28*16] = data_11_array[c23][d646][n646];
        end
    endgenerate
    generate 
        localparam integer d647 = 3;
        for (n647 = 0; n647 < 16; n647 = n647 + 1) 
        begin: outbit647
            assign data_11[n647 + d647*16 + c23*28*16] = data_11_array[c23][d647][n647];
        end
    endgenerate
    generate 
        localparam integer d648 = 4;
        for (n648 = 0; n648 < 16; n648 = n648 + 1) 
        begin: outbit648
            assign data_11[n648 + d648*16 + c23*28*16] = data_11_array[c23][d648][n648];
        end
    endgenerate
    generate 
        localparam integer d649 = 5;
        for (n649 = 0; n649 < 16; n649 = n649 + 1) 
        begin: outbit649
            assign data_11[n649 + d649*16 + c23*28*16] = data_11_array[c23][d649][n649];
        end
    endgenerate
    generate 
        localparam integer d650 = 6;
        for (n650 = 0; n650 < 16; n650 = n650 + 1) 
        begin: outbit650
            assign data_11[n650 + d650*16 + c23*28*16] = data_11_array[c23][d650][n650];
        end
    endgenerate
    generate 
        localparam integer d651 = 7;
        for (n651 = 0; n651 < 16; n651 = n651 + 1) 
        begin: outbit651
            assign data_11[n651 + d651*16 + c23*28*16] = data_11_array[c23][d651][n651];
        end
    endgenerate
    generate 
        localparam integer d652 = 8;
        for (n652 = 0; n652 < 16; n652 = n652 + 1) 
        begin: outbit652
            assign data_11[n652 + d652*16 + c23*28*16] = data_11_array[c23][d652][n652];
        end
    endgenerate
    generate 
        localparam integer d653 = 9;
        for (n653 = 0; n653 < 16; n653 = n653 + 1) 
        begin: outbit653
            assign data_11[n653 + d653*16 + c23*28*16] = data_11_array[c23][d653][n653];
        end
    endgenerate
    generate 
        localparam integer d654 = 10;
        for (n654 = 0; n654 < 16; n654 = n654 + 1) 
        begin: outbit654
            assign data_11[n654 + d654*16 + c23*28*16] = data_11_array[c23][d654][n654];
        end
    endgenerate
    generate 
        localparam integer d655 = 11;
        for (n655 = 0; n655 < 16; n655 = n655 + 1) 
        begin: outbit655
            assign data_11[n655 + d655*16 + c23*28*16] = data_11_array[c23][d655][n655];
        end
    endgenerate
    generate 
        localparam integer d656 = 12;
        for (n656 = 0; n656 < 16; n656 = n656 + 1) 
        begin: outbit656
            assign data_11[n656 + d656*16 + c23*28*16] = data_11_array[c23][d656][n656];
        end
    endgenerate
    generate 
        localparam integer d657 = 13;
        for (n657 = 0; n657 < 16; n657 = n657 + 1) 
        begin: outbit657
            assign data_11[n657 + d657*16 + c23*28*16] = data_11_array[c23][d657][n657];
        end
    endgenerate
    generate 
        localparam integer d658 = 14;
        for (n658 = 0; n658 < 16; n658 = n658 + 1) 
        begin: outbit658
            assign data_11[n658 + d658*16 + c23*28*16] = data_11_array[c23][d658][n658];
        end
    endgenerate
    generate 
        localparam integer d659 = 15;
        for (n659 = 0; n659 < 16; n659 = n659 + 1) 
        begin: outbit659
            assign data_11[n659 + d659*16 + c23*28*16] = data_11_array[c23][d659][n659];
        end
    endgenerate
    generate 
        localparam integer d660 = 16;
        for (n660 = 0; n660 < 16; n660 = n660 + 1) 
        begin: outbit660
            assign data_11[n660 + d660*16 + c23*28*16] = data_11_array[c23][d660][n660];
        end
    endgenerate
    generate 
        localparam integer d661 = 17;
        for (n661 = 0; n661 < 16; n661 = n661 + 1) 
        begin: outbit661
            assign data_11[n661 + d661*16 + c23*28*16] = data_11_array[c23][d661][n661];
        end
    endgenerate
    generate 
        localparam integer d662 = 18;
        for (n662 = 0; n662 < 16; n662 = n662 + 1) 
        begin: outbit662
            assign data_11[n662 + d662*16 + c23*28*16] = data_11_array[c23][d662][n662];
        end
    endgenerate
    generate 
        localparam integer d663 = 19;
        for (n663 = 0; n663 < 16; n663 = n663 + 1) 
        begin: outbit663
            assign data_11[n663 + d663*16 + c23*28*16] = data_11_array[c23][d663][n663];
        end
    endgenerate
    generate 
        localparam integer d664 = 20;
        for (n664 = 0; n664 < 16; n664 = n664 + 1) 
        begin: outbit664
            assign data_11[n664 + d664*16 + c23*28*16] = data_11_array[c23][d664][n664];
        end
    endgenerate
    generate 
        localparam integer d665 = 21;
        for (n665 = 0; n665 < 16; n665 = n665 + 1) 
        begin: outbit665
            assign data_11[n665 + d665*16 + c23*28*16] = data_11_array[c23][d665][n665];
        end
    endgenerate
    generate 
        localparam integer d666 = 22;
        for (n666 = 0; n666 < 16; n666 = n666 + 1) 
        begin: outbit666
            assign data_11[n666 + d666*16 + c23*28*16] = data_11_array[c23][d666][n666];
        end
    endgenerate
    generate 
        localparam integer d667 = 23;
        for (n667 = 0; n667 < 16; n667 = n667 + 1) 
        begin: outbit667
            assign data_11[n667 + d667*16 + c23*28*16] = data_11_array[c23][d667][n667];
        end
    endgenerate
    generate 
        localparam integer d668 = 24;
        for (n668 = 0; n668 < 16; n668 = n668 + 1) 
        begin: outbit668
            assign data_11[n668 + d668*16 + c23*28*16] = data_11_array[c23][d668][n668];
        end
    endgenerate
    generate 
        localparam integer d669 = 25;
        for (n669 = 0; n669 < 16; n669 = n669 + 1) 
        begin: outbit669
            assign data_11[n669 + d669*16 + c23*28*16] = data_11_array[c23][d669][n669];
        end
    endgenerate
    generate 
        localparam integer d670 = 26;
        for (n670 = 0; n670 < 16; n670 = n670 + 1) 
        begin: outbit670
            assign data_11[n670 + d670*16 + c23*28*16] = data_11_array[c23][d670][n670];
        end
    endgenerate
    generate 
        localparam integer d671 = 27;
        for (n671 = 0; n671 < 16; n671 = n671 + 1) 
        begin: outbit671
            assign data_11[n671 + d671*16 + c23*28*16] = data_11_array[c23][d671][n671];
        end
    endgenerate
    localparam integer c24 = 24;
    generate 
        localparam integer d672 = 0;
        for (n672 = 0; n672 < 16; n672 = n672 + 1) 
        begin: outbit672
            assign data_11[n672 + d672*16 + c24*28*16] = data_11_array[c24][d672][n672];
        end
    endgenerate
    generate 
        localparam integer d673 = 1;
        for (n673 = 0; n673 < 16; n673 = n673 + 1) 
        begin: outbit673
            assign data_11[n673 + d673*16 + c24*28*16] = data_11_array[c24][d673][n673];
        end
    endgenerate
    generate 
        localparam integer d674 = 2;
        for (n674 = 0; n674 < 16; n674 = n674 + 1) 
        begin: outbit674
            assign data_11[n674 + d674*16 + c24*28*16] = data_11_array[c24][d674][n674];
        end
    endgenerate
    generate 
        localparam integer d675 = 3;
        for (n675 = 0; n675 < 16; n675 = n675 + 1) 
        begin: outbit675
            assign data_11[n675 + d675*16 + c24*28*16] = data_11_array[c24][d675][n675];
        end
    endgenerate
    generate 
        localparam integer d676 = 4;
        for (n676 = 0; n676 < 16; n676 = n676 + 1) 
        begin: outbit676
            assign data_11[n676 + d676*16 + c24*28*16] = data_11_array[c24][d676][n676];
        end
    endgenerate
    generate 
        localparam integer d677 = 5;
        for (n677 = 0; n677 < 16; n677 = n677 + 1) 
        begin: outbit677
            assign data_11[n677 + d677*16 + c24*28*16] = data_11_array[c24][d677][n677];
        end
    endgenerate
    generate 
        localparam integer d678 = 6;
        for (n678 = 0; n678 < 16; n678 = n678 + 1) 
        begin: outbit678
            assign data_11[n678 + d678*16 + c24*28*16] = data_11_array[c24][d678][n678];
        end
    endgenerate
    generate 
        localparam integer d679 = 7;
        for (n679 = 0; n679 < 16; n679 = n679 + 1) 
        begin: outbit679
            assign data_11[n679 + d679*16 + c24*28*16] = data_11_array[c24][d679][n679];
        end
    endgenerate
    generate 
        localparam integer d680 = 8;
        for (n680 = 0; n680 < 16; n680 = n680 + 1) 
        begin: outbit680
            assign data_11[n680 + d680*16 + c24*28*16] = data_11_array[c24][d680][n680];
        end
    endgenerate
    generate 
        localparam integer d681 = 9;
        for (n681 = 0; n681 < 16; n681 = n681 + 1) 
        begin: outbit681
            assign data_11[n681 + d681*16 + c24*28*16] = data_11_array[c24][d681][n681];
        end
    endgenerate
    generate 
        localparam integer d682 = 10;
        for (n682 = 0; n682 < 16; n682 = n682 + 1) 
        begin: outbit682
            assign data_11[n682 + d682*16 + c24*28*16] = data_11_array[c24][d682][n682];
        end
    endgenerate
    generate 
        localparam integer d683 = 11;
        for (n683 = 0; n683 < 16; n683 = n683 + 1) 
        begin: outbit683
            assign data_11[n683 + d683*16 + c24*28*16] = data_11_array[c24][d683][n683];
        end
    endgenerate
    generate 
        localparam integer d684 = 12;
        for (n684 = 0; n684 < 16; n684 = n684 + 1) 
        begin: outbit684
            assign data_11[n684 + d684*16 + c24*28*16] = data_11_array[c24][d684][n684];
        end
    endgenerate
    generate 
        localparam integer d685 = 13;
        for (n685 = 0; n685 < 16; n685 = n685 + 1) 
        begin: outbit685
            assign data_11[n685 + d685*16 + c24*28*16] = data_11_array[c24][d685][n685];
        end
    endgenerate
    generate 
        localparam integer d686 = 14;
        for (n686 = 0; n686 < 16; n686 = n686 + 1) 
        begin: outbit686
            assign data_11[n686 + d686*16 + c24*28*16] = data_11_array[c24][d686][n686];
        end
    endgenerate
    generate 
        localparam integer d687 = 15;
        for (n687 = 0; n687 < 16; n687 = n687 + 1) 
        begin: outbit687
            assign data_11[n687 + d687*16 + c24*28*16] = data_11_array[c24][d687][n687];
        end
    endgenerate
    generate 
        localparam integer d688 = 16;
        for (n688 = 0; n688 < 16; n688 = n688 + 1) 
        begin: outbit688
            assign data_11[n688 + d688*16 + c24*28*16] = data_11_array[c24][d688][n688];
        end
    endgenerate
    generate 
        localparam integer d689 = 17;
        for (n689 = 0; n689 < 16; n689 = n689 + 1) 
        begin: outbit689
            assign data_11[n689 + d689*16 + c24*28*16] = data_11_array[c24][d689][n689];
        end
    endgenerate
    generate 
        localparam integer d690 = 18;
        for (n690 = 0; n690 < 16; n690 = n690 + 1) 
        begin: outbit690
            assign data_11[n690 + d690*16 + c24*28*16] = data_11_array[c24][d690][n690];
        end
    endgenerate
    generate 
        localparam integer d691 = 19;
        for (n691 = 0; n691 < 16; n691 = n691 + 1) 
        begin: outbit691
            assign data_11[n691 + d691*16 + c24*28*16] = data_11_array[c24][d691][n691];
        end
    endgenerate
    generate 
        localparam integer d692 = 20;
        for (n692 = 0; n692 < 16; n692 = n692 + 1) 
        begin: outbit692
            assign data_11[n692 + d692*16 + c24*28*16] = data_11_array[c24][d692][n692];
        end
    endgenerate
    generate 
        localparam integer d693 = 21;
        for (n693 = 0; n693 < 16; n693 = n693 + 1) 
        begin: outbit693
            assign data_11[n693 + d693*16 + c24*28*16] = data_11_array[c24][d693][n693];
        end
    endgenerate
    generate 
        localparam integer d694 = 22;
        for (n694 = 0; n694 < 16; n694 = n694 + 1) 
        begin: outbit694
            assign data_11[n694 + d694*16 + c24*28*16] = data_11_array[c24][d694][n694];
        end
    endgenerate
    generate 
        localparam integer d695 = 23;
        for (n695 = 0; n695 < 16; n695 = n695 + 1) 
        begin: outbit695
            assign data_11[n695 + d695*16 + c24*28*16] = data_11_array[c24][d695][n695];
        end
    endgenerate
    generate 
        localparam integer d696 = 24;
        for (n696 = 0; n696 < 16; n696 = n696 + 1) 
        begin: outbit696
            assign data_11[n696 + d696*16 + c24*28*16] = data_11_array[c24][d696][n696];
        end
    endgenerate
    generate 
        localparam integer d697 = 25;
        for (n697 = 0; n697 < 16; n697 = n697 + 1) 
        begin: outbit697
            assign data_11[n697 + d697*16 + c24*28*16] = data_11_array[c24][d697][n697];
        end
    endgenerate
    generate 
        localparam integer d698 = 26;
        for (n698 = 0; n698 < 16; n698 = n698 + 1) 
        begin: outbit698
            assign data_11[n698 + d698*16 + c24*28*16] = data_11_array[c24][d698][n698];
        end
    endgenerate
    generate 
        localparam integer d699 = 27;
        for (n699 = 0; n699 < 16; n699 = n699 + 1) 
        begin: outbit699
            assign data_11[n699 + d699*16 + c24*28*16] = data_11_array[c24][d699][n699];
        end
    endgenerate
    localparam integer c25 = 25;
    generate 
        localparam integer d700 = 0;
        for (n700 = 0; n700 < 16; n700 = n700 + 1) 
        begin: outbit700
            assign data_11[n700 + d700*16 + c25*28*16] = data_11_array[c25][d700][n700];
        end
    endgenerate
    generate 
        localparam integer d701 = 1;
        for (n701 = 0; n701 < 16; n701 = n701 + 1) 
        begin: outbit701
            assign data_11[n701 + d701*16 + c25*28*16] = data_11_array[c25][d701][n701];
        end
    endgenerate
    generate 
        localparam integer d702 = 2;
        for (n702 = 0; n702 < 16; n702 = n702 + 1) 
        begin: outbit702
            assign data_11[n702 + d702*16 + c25*28*16] = data_11_array[c25][d702][n702];
        end
    endgenerate
    generate 
        localparam integer d703 = 3;
        for (n703 = 0; n703 < 16; n703 = n703 + 1) 
        begin: outbit703
            assign data_11[n703 + d703*16 + c25*28*16] = data_11_array[c25][d703][n703];
        end
    endgenerate
    generate 
        localparam integer d704 = 4;
        for (n704 = 0; n704 < 16; n704 = n704 + 1) 
        begin: outbit704
            assign data_11[n704 + d704*16 + c25*28*16] = data_11_array[c25][d704][n704];
        end
    endgenerate
    generate 
        localparam integer d705 = 5;
        for (n705 = 0; n705 < 16; n705 = n705 + 1) 
        begin: outbit705
            assign data_11[n705 + d705*16 + c25*28*16] = data_11_array[c25][d705][n705];
        end
    endgenerate
    generate 
        localparam integer d706 = 6;
        for (n706 = 0; n706 < 16; n706 = n706 + 1) 
        begin: outbit706
            assign data_11[n706 + d706*16 + c25*28*16] = data_11_array[c25][d706][n706];
        end
    endgenerate
    generate 
        localparam integer d707 = 7;
        for (n707 = 0; n707 < 16; n707 = n707 + 1) 
        begin: outbit707
            assign data_11[n707 + d707*16 + c25*28*16] = data_11_array[c25][d707][n707];
        end
    endgenerate
    generate 
        localparam integer d708 = 8;
        for (n708 = 0; n708 < 16; n708 = n708 + 1) 
        begin: outbit708
            assign data_11[n708 + d708*16 + c25*28*16] = data_11_array[c25][d708][n708];
        end
    endgenerate
    generate 
        localparam integer d709 = 9;
        for (n709 = 0; n709 < 16; n709 = n709 + 1) 
        begin: outbit709
            assign data_11[n709 + d709*16 + c25*28*16] = data_11_array[c25][d709][n709];
        end
    endgenerate
    generate 
        localparam integer d710 = 10;
        for (n710 = 0; n710 < 16; n710 = n710 + 1) 
        begin: outbit710
            assign data_11[n710 + d710*16 + c25*28*16] = data_11_array[c25][d710][n710];
        end
    endgenerate
    generate 
        localparam integer d711 = 11;
        for (n711 = 0; n711 < 16; n711 = n711 + 1) 
        begin: outbit711
            assign data_11[n711 + d711*16 + c25*28*16] = data_11_array[c25][d711][n711];
        end
    endgenerate
    generate 
        localparam integer d712 = 12;
        for (n712 = 0; n712 < 16; n712 = n712 + 1) 
        begin: outbit712
            assign data_11[n712 + d712*16 + c25*28*16] = data_11_array[c25][d712][n712];
        end
    endgenerate
    generate 
        localparam integer d713 = 13;
        for (n713 = 0; n713 < 16; n713 = n713 + 1) 
        begin: outbit713
            assign data_11[n713 + d713*16 + c25*28*16] = data_11_array[c25][d713][n713];
        end
    endgenerate
    generate 
        localparam integer d714 = 14;
        for (n714 = 0; n714 < 16; n714 = n714 + 1) 
        begin: outbit714
            assign data_11[n714 + d714*16 + c25*28*16] = data_11_array[c25][d714][n714];
        end
    endgenerate
    generate 
        localparam integer d715 = 15;
        for (n715 = 0; n715 < 16; n715 = n715 + 1) 
        begin: outbit715
            assign data_11[n715 + d715*16 + c25*28*16] = data_11_array[c25][d715][n715];
        end
    endgenerate
    generate 
        localparam integer d716 = 16;
        for (n716 = 0; n716 < 16; n716 = n716 + 1) 
        begin: outbit716
            assign data_11[n716 + d716*16 + c25*28*16] = data_11_array[c25][d716][n716];
        end
    endgenerate
    generate 
        localparam integer d717 = 17;
        for (n717 = 0; n717 < 16; n717 = n717 + 1) 
        begin: outbit717
            assign data_11[n717 + d717*16 + c25*28*16] = data_11_array[c25][d717][n717];
        end
    endgenerate
    generate 
        localparam integer d718 = 18;
        for (n718 = 0; n718 < 16; n718 = n718 + 1) 
        begin: outbit718
            assign data_11[n718 + d718*16 + c25*28*16] = data_11_array[c25][d718][n718];
        end
    endgenerate
    generate 
        localparam integer d719 = 19;
        for (n719 = 0; n719 < 16; n719 = n719 + 1) 
        begin: outbit719
            assign data_11[n719 + d719*16 + c25*28*16] = data_11_array[c25][d719][n719];
        end
    endgenerate
    generate 
        localparam integer d720 = 20;
        for (n720 = 0; n720 < 16; n720 = n720 + 1) 
        begin: outbit720
            assign data_11[n720 + d720*16 + c25*28*16] = data_11_array[c25][d720][n720];
        end
    endgenerate
    generate 
        localparam integer d721 = 21;
        for (n721 = 0; n721 < 16; n721 = n721 + 1) 
        begin: outbit721
            assign data_11[n721 + d721*16 + c25*28*16] = data_11_array[c25][d721][n721];
        end
    endgenerate
    generate 
        localparam integer d722 = 22;
        for (n722 = 0; n722 < 16; n722 = n722 + 1) 
        begin: outbit722
            assign data_11[n722 + d722*16 + c25*28*16] = data_11_array[c25][d722][n722];
        end
    endgenerate
    generate 
        localparam integer d723 = 23;
        for (n723 = 0; n723 < 16; n723 = n723 + 1) 
        begin: outbit723
            assign data_11[n723 + d723*16 + c25*28*16] = data_11_array[c25][d723][n723];
        end
    endgenerate
    generate 
        localparam integer d724 = 24;
        for (n724 = 0; n724 < 16; n724 = n724 + 1) 
        begin: outbit724
            assign data_11[n724 + d724*16 + c25*28*16] = data_11_array[c25][d724][n724];
        end
    endgenerate
    generate 
        localparam integer d725 = 25;
        for (n725 = 0; n725 < 16; n725 = n725 + 1) 
        begin: outbit725
            assign data_11[n725 + d725*16 + c25*28*16] = data_11_array[c25][d725][n725];
        end
    endgenerate
    generate 
        localparam integer d726 = 26;
        for (n726 = 0; n726 < 16; n726 = n726 + 1) 
        begin: outbit726
            assign data_11[n726 + d726*16 + c25*28*16] = data_11_array[c25][d726][n726];
        end
    endgenerate
    generate 
        localparam integer d727 = 27;
        for (n727 = 0; n727 < 16; n727 = n727 + 1) 
        begin: outbit727
            assign data_11[n727 + d727*16 + c25*28*16] = data_11_array[c25][d727][n727];
        end
    endgenerate
    localparam integer c26 = 26;
    generate 
        localparam integer d728 = 0;
        for (n728 = 0; n728 < 16; n728 = n728 + 1) 
        begin: outbit728
            assign data_11[n728 + d728*16 + c26*28*16] = data_11_array[c26][d728][n728];
        end
    endgenerate
    generate 
        localparam integer d729 = 1;
        for (n729 = 0; n729 < 16; n729 = n729 + 1) 
        begin: outbit729
            assign data_11[n729 + d729*16 + c26*28*16] = data_11_array[c26][d729][n729];
        end
    endgenerate
    generate 
        localparam integer d730 = 2;
        for (n730 = 0; n730 < 16; n730 = n730 + 1) 
        begin: outbit730
            assign data_11[n730 + d730*16 + c26*28*16] = data_11_array[c26][d730][n730];
        end
    endgenerate
    generate 
        localparam integer d731 = 3;
        for (n731 = 0; n731 < 16; n731 = n731 + 1) 
        begin: outbit731
            assign data_11[n731 + d731*16 + c26*28*16] = data_11_array[c26][d731][n731];
        end
    endgenerate
    generate 
        localparam integer d732 = 4;
        for (n732 = 0; n732 < 16; n732 = n732 + 1) 
        begin: outbit732
            assign data_11[n732 + d732*16 + c26*28*16] = data_11_array[c26][d732][n732];
        end
    endgenerate
    generate 
        localparam integer d733 = 5;
        for (n733 = 0; n733 < 16; n733 = n733 + 1) 
        begin: outbit733
            assign data_11[n733 + d733*16 + c26*28*16] = data_11_array[c26][d733][n733];
        end
    endgenerate
    generate 
        localparam integer d734 = 6;
        for (n734 = 0; n734 < 16; n734 = n734 + 1) 
        begin: outbit734
            assign data_11[n734 + d734*16 + c26*28*16] = data_11_array[c26][d734][n734];
        end
    endgenerate
    generate 
        localparam integer d735 = 7;
        for (n735 = 0; n735 < 16; n735 = n735 + 1) 
        begin: outbit735
            assign data_11[n735 + d735*16 + c26*28*16] = data_11_array[c26][d735][n735];
        end
    endgenerate
    generate 
        localparam integer d736 = 8;
        for (n736 = 0; n736 < 16; n736 = n736 + 1) 
        begin: outbit736
            assign data_11[n736 + d736*16 + c26*28*16] = data_11_array[c26][d736][n736];
        end
    endgenerate
    generate 
        localparam integer d737 = 9;
        for (n737 = 0; n737 < 16; n737 = n737 + 1) 
        begin: outbit737
            assign data_11[n737 + d737*16 + c26*28*16] = data_11_array[c26][d737][n737];
        end
    endgenerate
    generate 
        localparam integer d738 = 10;
        for (n738 = 0; n738 < 16; n738 = n738 + 1) 
        begin: outbit738
            assign data_11[n738 + d738*16 + c26*28*16] = data_11_array[c26][d738][n738];
        end
    endgenerate
    generate 
        localparam integer d739 = 11;
        for (n739 = 0; n739 < 16; n739 = n739 + 1) 
        begin: outbit739
            assign data_11[n739 + d739*16 + c26*28*16] = data_11_array[c26][d739][n739];
        end
    endgenerate
    generate 
        localparam integer d740 = 12;
        for (n740 = 0; n740 < 16; n740 = n740 + 1) 
        begin: outbit740
            assign data_11[n740 + d740*16 + c26*28*16] = data_11_array[c26][d740][n740];
        end
    endgenerate
    generate 
        localparam integer d741 = 13;
        for (n741 = 0; n741 < 16; n741 = n741 + 1) 
        begin: outbit741
            assign data_11[n741 + d741*16 + c26*28*16] = data_11_array[c26][d741][n741];
        end
    endgenerate
    generate 
        localparam integer d742 = 14;
        for (n742 = 0; n742 < 16; n742 = n742 + 1) 
        begin: outbit742
            assign data_11[n742 + d742*16 + c26*28*16] = data_11_array[c26][d742][n742];
        end
    endgenerate
    generate 
        localparam integer d743 = 15;
        for (n743 = 0; n743 < 16; n743 = n743 + 1) 
        begin: outbit743
            assign data_11[n743 + d743*16 + c26*28*16] = data_11_array[c26][d743][n743];
        end
    endgenerate
    generate 
        localparam integer d744 = 16;
        for (n744 = 0; n744 < 16; n744 = n744 + 1) 
        begin: outbit744
            assign data_11[n744 + d744*16 + c26*28*16] = data_11_array[c26][d744][n744];
        end
    endgenerate
    generate 
        localparam integer d745 = 17;
        for (n745 = 0; n745 < 16; n745 = n745 + 1) 
        begin: outbit745
            assign data_11[n745 + d745*16 + c26*28*16] = data_11_array[c26][d745][n745];
        end
    endgenerate
    generate 
        localparam integer d746 = 18;
        for (n746 = 0; n746 < 16; n746 = n746 + 1) 
        begin: outbit746
            assign data_11[n746 + d746*16 + c26*28*16] = data_11_array[c26][d746][n746];
        end
    endgenerate
    generate 
        localparam integer d747 = 19;
        for (n747 = 0; n747 < 16; n747 = n747 + 1) 
        begin: outbit747
            assign data_11[n747 + d747*16 + c26*28*16] = data_11_array[c26][d747][n747];
        end
    endgenerate
    generate 
        localparam integer d748 = 20;
        for (n748 = 0; n748 < 16; n748 = n748 + 1) 
        begin: outbit748
            assign data_11[n748 + d748*16 + c26*28*16] = data_11_array[c26][d748][n748];
        end
    endgenerate
    generate 
        localparam integer d749 = 21;
        for (n749 = 0; n749 < 16; n749 = n749 + 1) 
        begin: outbit749
            assign data_11[n749 + d749*16 + c26*28*16] = data_11_array[c26][d749][n749];
        end
    endgenerate
    generate 
        localparam integer d750 = 22;
        for (n750 = 0; n750 < 16; n750 = n750 + 1) 
        begin: outbit750
            assign data_11[n750 + d750*16 + c26*28*16] = data_11_array[c26][d750][n750];
        end
    endgenerate
    generate 
        localparam integer d751 = 23;
        for (n751 = 0; n751 < 16; n751 = n751 + 1) 
        begin: outbit751
            assign data_11[n751 + d751*16 + c26*28*16] = data_11_array[c26][d751][n751];
        end
    endgenerate
    generate 
        localparam integer d752 = 24;
        for (n752 = 0; n752 < 16; n752 = n752 + 1) 
        begin: outbit752
            assign data_11[n752 + d752*16 + c26*28*16] = data_11_array[c26][d752][n752];
        end
    endgenerate
    generate 
        localparam integer d753 = 25;
        for (n753 = 0; n753 < 16; n753 = n753 + 1) 
        begin: outbit753
            assign data_11[n753 + d753*16 + c26*28*16] = data_11_array[c26][d753][n753];
        end
    endgenerate
    generate 
        localparam integer d754 = 26;
        for (n754 = 0; n754 < 16; n754 = n754 + 1) 
        begin: outbit754
            assign data_11[n754 + d754*16 + c26*28*16] = data_11_array[c26][d754][n754];
        end
    endgenerate
    generate 
        localparam integer d755 = 27;
        for (n755 = 0; n755 < 16; n755 = n755 + 1) 
        begin: outbit755
            assign data_11[n755 + d755*16 + c26*28*16] = data_11_array[c26][d755][n755];
        end
    endgenerate
    localparam integer c27 = 27;
    generate 
        localparam integer d756 = 0;
        for (n756 = 0; n756 < 16; n756 = n756 + 1) 
        begin: outbit756
            assign data_11[n756 + d756*16 + c27*28*16] = data_11_array[c27][d756][n756];
        end
    endgenerate
    generate 
        localparam integer d757 = 1;
        for (n757 = 0; n757 < 16; n757 = n757 + 1) 
        begin: outbit757
            assign data_11[n757 + d757*16 + c27*28*16] = data_11_array[c27][d757][n757];
        end
    endgenerate
    generate 
        localparam integer d758 = 2;
        for (n758 = 0; n758 < 16; n758 = n758 + 1) 
        begin: outbit758
            assign data_11[n758 + d758*16 + c27*28*16] = data_11_array[c27][d758][n758];
        end
    endgenerate
    generate 
        localparam integer d759 = 3;
        for (n759 = 0; n759 < 16; n759 = n759 + 1) 
        begin: outbit759
            assign data_11[n759 + d759*16 + c27*28*16] = data_11_array[c27][d759][n759];
        end
    endgenerate
    generate 
        localparam integer d760 = 4;
        for (n760 = 0; n760 < 16; n760 = n760 + 1) 
        begin: outbit760
            assign data_11[n760 + d760*16 + c27*28*16] = data_11_array[c27][d760][n760];
        end
    endgenerate
    generate 
        localparam integer d761 = 5;
        for (n761 = 0; n761 < 16; n761 = n761 + 1) 
        begin: outbit761
            assign data_11[n761 + d761*16 + c27*28*16] = data_11_array[c27][d761][n761];
        end
    endgenerate
    generate 
        localparam integer d762 = 6;
        for (n762 = 0; n762 < 16; n762 = n762 + 1) 
        begin: outbit762
            assign data_11[n762 + d762*16 + c27*28*16] = data_11_array[c27][d762][n762];
        end
    endgenerate
    generate 
        localparam integer d763 = 7;
        for (n763 = 0; n763 < 16; n763 = n763 + 1) 
        begin: outbit763
            assign data_11[n763 + d763*16 + c27*28*16] = data_11_array[c27][d763][n763];
        end
    endgenerate
    generate 
        localparam integer d764 = 8;
        for (n764 = 0; n764 < 16; n764 = n764 + 1) 
        begin: outbit764
            assign data_11[n764 + d764*16 + c27*28*16] = data_11_array[c27][d764][n764];
        end
    endgenerate
    generate 
        localparam integer d765 = 9;
        for (n765 = 0; n765 < 16; n765 = n765 + 1) 
        begin: outbit765
            assign data_11[n765 + d765*16 + c27*28*16] = data_11_array[c27][d765][n765];
        end
    endgenerate
    generate 
        localparam integer d766 = 10;
        for (n766 = 0; n766 < 16; n766 = n766 + 1) 
        begin: outbit766
            assign data_11[n766 + d766*16 + c27*28*16] = data_11_array[c27][d766][n766];
        end
    endgenerate
    generate 
        localparam integer d767 = 11;
        for (n767 = 0; n767 < 16; n767 = n767 + 1) 
        begin: outbit767
            assign data_11[n767 + d767*16 + c27*28*16] = data_11_array[c27][d767][n767];
        end
    endgenerate
    generate 
        localparam integer d768 = 12;
        for (n768 = 0; n768 < 16; n768 = n768 + 1) 
        begin: outbit768
            assign data_11[n768 + d768*16 + c27*28*16] = data_11_array[c27][d768][n768];
        end
    endgenerate
    generate 
        localparam integer d769 = 13;
        for (n769 = 0; n769 < 16; n769 = n769 + 1) 
        begin: outbit769
            assign data_11[n769 + d769*16 + c27*28*16] = data_11_array[c27][d769][n769];
        end
    endgenerate
    generate 
        localparam integer d770 = 14;
        for (n770 = 0; n770 < 16; n770 = n770 + 1) 
        begin: outbit770
            assign data_11[n770 + d770*16 + c27*28*16] = data_11_array[c27][d770][n770];
        end
    endgenerate
    generate 
        localparam integer d771 = 15;
        for (n771 = 0; n771 < 16; n771 = n771 + 1) 
        begin: outbit771
            assign data_11[n771 + d771*16 + c27*28*16] = data_11_array[c27][d771][n771];
        end
    endgenerate
    generate 
        localparam integer d772 = 16;
        for (n772 = 0; n772 < 16; n772 = n772 + 1) 
        begin: outbit772
            assign data_11[n772 + d772*16 + c27*28*16] = data_11_array[c27][d772][n772];
        end
    endgenerate
    generate 
        localparam integer d773 = 17;
        for (n773 = 0; n773 < 16; n773 = n773 + 1) 
        begin: outbit773
            assign data_11[n773 + d773*16 + c27*28*16] = data_11_array[c27][d773][n773];
        end
    endgenerate
    generate 
        localparam integer d774 = 18;
        for (n774 = 0; n774 < 16; n774 = n774 + 1) 
        begin: outbit774
            assign data_11[n774 + d774*16 + c27*28*16] = data_11_array[c27][d774][n774];
        end
    endgenerate
    generate 
        localparam integer d775 = 19;
        for (n775 = 0; n775 < 16; n775 = n775 + 1) 
        begin: outbit775
            assign data_11[n775 + d775*16 + c27*28*16] = data_11_array[c27][d775][n775];
        end
    endgenerate
    generate 
        localparam integer d776 = 20;
        for (n776 = 0; n776 < 16; n776 = n776 + 1) 
        begin: outbit776
            assign data_11[n776 + d776*16 + c27*28*16] = data_11_array[c27][d776][n776];
        end
    endgenerate
    generate 
        localparam integer d777 = 21;
        for (n777 = 0; n777 < 16; n777 = n777 + 1) 
        begin: outbit777
            assign data_11[n777 + d777*16 + c27*28*16] = data_11_array[c27][d777][n777];
        end
    endgenerate
    generate 
        localparam integer d778 = 22;
        for (n778 = 0; n778 < 16; n778 = n778 + 1) 
        begin: outbit778
            assign data_11[n778 + d778*16 + c27*28*16] = data_11_array[c27][d778][n778];
        end
    endgenerate
    generate 
        localparam integer d779 = 23;
        for (n779 = 0; n779 < 16; n779 = n779 + 1) 
        begin: outbit779
            assign data_11[n779 + d779*16 + c27*28*16] = data_11_array[c27][d779][n779];
        end
    endgenerate
    generate 
        localparam integer d780 = 24;
        for (n780 = 0; n780 < 16; n780 = n780 + 1) 
        begin: outbit780
            assign data_11[n780 + d780*16 + c27*28*16] = data_11_array[c27][d780][n780];
        end
    endgenerate
    generate 
        localparam integer d781 = 25;
        for (n781 = 0; n781 < 16; n781 = n781 + 1) 
        begin: outbit781
            assign data_11[n781 + d781*16 + c27*28*16] = data_11_array[c27][d781][n781];
        end
    endgenerate
    generate 
        localparam integer d782 = 26;
        for (n782 = 0; n782 < 16; n782 = n782 + 1) 
        begin: outbit782
            assign data_11[n782 + d782*16 + c27*28*16] = data_11_array[c27][d782][n782];
        end
    endgenerate
    generate 
        localparam integer d783 = 27;
        for (n783 = 0; n783 < 16; n783 = n783 + 1) 
        begin: outbit783
            assign data_11[n783 + d783*16 + c27*28*16] = data_11_array[c27][d783][n783];
        end
    endgenerate

endmodule

////CONVOLUTION LAYER 1 | FEATURE MAP 4
module Conv1_feature4 (
    data,
    feature4Weight_0,
    feature4Weight_1,
    feature4Weight_2,
    feature4Weight_3,
    feature4Weight_4,
    feature4Weight_5,
    feature4Weight_6,
    feature4Weight_7,
    feature4Weight_8,
    feature4Weight_9,
    feature4Weight_10,
    feature4Weight_11,
    feature4Weight_12,
    feature4Weight_13,
    feature4Weight_14,
    feature4Weight_15,
    feature4Weight_16,
    feature4Weight_17,
    feature4Weight_18,
    feature4Weight_19,
    feature4Weight_20,
    feature4Weight_21,
    feature4Weight_22,
    feature4Weight_23,
    feature4Weight_24,
    feature4Bias,
    data_11);

  parameter TEST_DATA = 784*16,
    FP_LENGTH = 16;
  input [TEST_DATA - 1:0] data;
  input [FP_LENGTH - 1:0] feature4Weight_0, feature4Weight_1, feature4Weight_2, feature4Weight_3, feature4Weight_4, feature4Weight_5, feature4Weight_6, feature4Weight_7, feature4Weight_8, feature4Weight_9, feature4Weight_10, feature4Weight_11, feature4Weight_12, feature4Weight_13, feature4Weight_14, feature4Weight_15, feature4Weight_16, feature4Weight_17, feature4Weight_18, feature4Weight_19, feature4Weight_20, feature4Weight_21, feature4Weight_22, feature4Weight_23, feature4Weight_24, feature4Bias;
  output [576*16 - 1:0] data_11;    
  
  wire [FP_LENGTH - 1:0] data_array [0:27][0:27];
  wire [FP_LENGTH - 1:0] data_11_array [0:23][0:23];
  wire [FP_LENGTH - 1:0] multi0 [0:24][0:23], multi1 [0:24][0:23], multi2 [0:24][0:23], multi3 [0:24][0:23], multi4 [0:24][0:23], multi5 [0:24][0:23], multi6 [0:24][0:23], multi7 [0:24][0:23], multi8 [0:24][0:23], multi9 [0:24][0:23], multi10 [0:24][0:23], multi11 [0:24][0:23], multi12 [0:24][0:23], multi13 [0:24][0:23], multi14 [0:24][0:23], multi15 [0:24][0:23], multi16 [0:24][0:23], multi17 [0:24][0:23], multi18 [0:24][0:23], multi19 [0:24][0:23], multi20 [0:24][0:23], multi21 [0:24][0:23], multi22 [0:24][0:23], multi23 [0:24][0:23], multi24 [0:24][0:23];
  wire [FP_LENGTH - 1:0] sum0 [0:23][0:23], sum1 [0:23][0:23], sum2 [0:23][0:23], sum3 [0:23][0:23], sum4 [0:23][0:23], sum5 [0:23][0:23], sum6 [0:23][0:23], sum7 [0:23][0:23], sum8 [0:23][0:23], sum9 [0:23][0:23], sum10 [0:23][0:23], sum11 [0:23][0:23], sum12 [0:23][0:23], sum13 [0:23][0:23], sum14 [0:23][0:23], sum15 [0:23][0:23], sum16 [0:23][0:23], sum17 [0:23][0:23], sum18 [0:23][0:23], sum19 [0:23][0:23], sum20 [0:23][0:23], sum21 [0:23][0:23], sum22 [0:23][0:23], sum23 [0:23][0:23], sum24 [0:23][0:23];
//  integer a, b, c; ///a = ROW, b = COLUMN, c = 16 bit Value
  
//  initial begin
//    for (a = 0; a < 28; a = a + 1) begin
//        for (b = 0; b < 28; b = b + 1) begin
//            for (c = 15; c >= 0; c = c - 1) begin
//                data_array[a][b][c] = data[c + b*16 + a*28*16];
//            end
//        end
//    end
    
//    forever begin
//        for (a = 0; a < 28; a = a + 1) begin
//            for (b = 0; b < 28; b = b + 1) begin
//                for (c = 15; c >= 0; c = c - 1) begin
//                   data_11[c + b*16 + a*28*16] = data_11_array[a][b][c];
//                end
//            end
//        end
//    end
//  end
  
  
  
  genvar i0, i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20, i21, i22, i23, m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15,m16,m17,m18,m19,m20,m21,m22,m23,m24,m25,m26,m27,m28,m29,m30,m31,m32,m33,m34,m35,m36,m37,m38,m39,m40,m41,m42,m43,m44,m45,m46,m47,m48,m49,m50,m51,m52,m53,m54,m55,m56,m57,m58,m59,m60,m61,m62,m63,m64,m65,m66,m67,m68,m69,m70,m71,m72,m73,m74,m75,m76,m77,m78,m79,m80,m81,m82,m83,m84,m85,m86,m87,m88,m89,m90,m91,m92,m93,m94,m95,m96,m97,m98,m99,m100,m101,m102,m103,m104,m105,m106,m107,m108,m109,m110,m111,m112,m113,m114,m115,m116,m117,m118,m119,m120,m121,m122,m123,m124,m125,m126,m127,m128,m129,m130,m131,m132,m133,m134,m135,m136,m137,m138,m139,m140,m141,m142,m143,m144,m145,m146,m147,m148,m149,m150,m151,m152,m153,m154,m155,m156,m157,m158,m159,m160,m161,m162,m163,m164,m165,m166,m167,m168,m169,m170,m171,m172,m173,m174,m175,m176,m177,m178,m179,m180,m181,m182,m183,m184,m185,m186,m187,m188,m189,m190,m191,m192,m193,m194,m195,m196,m197,m198,m199,m200,m201,m202,m203,m204,m205,m206,m207,m208,m209,m210,m211,m212,m213,m214,m215,m216,m217,m218,m219,m220,m221,m222,m223,m224,m225,m226,m227,m228,m229,m230,m231,m232,m233,m234,m235,m236,m237,m238,m239,m240,m241,m242,m243,m244,m245,m246,m247,m248,m249,m250,m251,m252,m253,m254,m255,m256,m257,m258,m259,m260,m261,m262,m263,m264,m265,m266,m267,m268,m269,m270,m271,m272,m273,m274,m275,m276,m277,m278,m279,m280,m281,m282,m283,m284,m285,m286,m287,m288,m289,m290,m291,m292,m293,m294,m295,m296,m297,m298,m299,m300,m301,m302,m303,m304,m305,m306,m307,m308,m309,m310,m311,m312,m313,m314,m315,m316,m317,m318,m319,m320,m321,m322,m323,m324,m325,m326,m327,m328,m329,m330,m331,m332,m333,m334,m335,m336,m337,m338,m339,m340,m341,m342,m343,m344,m345,m346,m347,m348,m349,m350,m351,m352,m353,m354,m355,m356,m357,m358,m359,m360,m361,m362,m363,m364,m365,m366,m367,m368,m369,m370,m371,m372,m373,m374,m375,m376,m377,m378,m379,m380,m381,m382,m383,m384,m385,m386,m387,m388,m389,m390,m391,m392,m393,m394,m395,m396,m397,m398,m399,m400,m401,m402,m403,m404,m405,m406,m407,m408,m409,m410,m411,m412,m413,m414,m415,m416,m417,m418,m419,m420,m421,m422,m423,m424,m425,m426,m427,m428,m429,m430,m431,m432,m433,m434,m435,m436,m437,m438,m439,m440,m441,m442,m443,m444,m445,m446,m447,m448,m449,m450,m451,m452,m453,m454,m455,m456,m457,m458,m459,m460,m461,m462,m463,m464,m465,m466,m467,m468,m469,m470,m471,m472,m473,m474,m475,m476,m477,m478,m479,m480,m481,m482,m483,m484,m485,m486,m487,m488,m489,m490,m491,m492,m493,m494,m495,m496,m497,m498,m499,m500,m501,m502,m503,m504,m505,m506,m507,m508,m509,m510,m511,m512,m513,m514,m515,m516,m517,m518,m519,m520,m521,m522,m523,m524,m525,m526,m527,m528,m529,m530,m531,m532,m533,m534,m535,m536,m537,m538,m539,m540,m541,m542,m543,m544,m545,m546,m547,m548,m549,m550,m551,m552,m553,m554,m555,m556,m557,m558,m559,m560,m561,m562,m563,m564,m565,m566,m567,m568,m569,m570,m571,m572,m573,m574,m575,m576,m577,m578,m579,m580,m581,m582,m583,m584,m585,m586,m587,m588,m589,m590,m591,m592,m593,m594,m595,m596,m597,m598,m599,m600,m601,m602,m603,m604,m605,m606,m607,m608,m609,m610,m611,m612,m613,m614,m615,m616,m617,m618,m619,m620,m621,m622,m623,m624,m625,m626,m627,m628,m629,m630,m631,m632,m633,m634,m635,m636,m637,m638,m639,m640,m641,m642,m643,m644,m645,m646,m647,m648,m649,m650,m651,m652,m653,m654,m655,m656,m657,m658,m659,m660,m661,m662,m663,m664,m665,m666,m667,m668,m669,m670,m671,m672,m673,m674,m675,m676,m677,m678,m679,m680,m681,m682,m683,m684,m685,m686,m687,m688,m689,m690,m691,m692,m693,m694,m695,m696,m697,m698,m699,m700,m701,m702,m703,m704,m705,m706,m707,m708,m709,m710,m711,m712,m713,m714,m715,m716,m717,m718,m719,m720,m721,m722,m723,m724,m725,m726,m727,m728,m729,m730,m731,m732,m733,m734,m735,m736,m737,m738,m739,m740,m741,m742,m743,m744,m745,m746,m747,m748,m749,m750,m751,m752,m753,m754,m755,m756,m757,m758,m759,m760,m761,m762,m763,m764,m765,m766,m767,m768,m769,m770,m771,m772,m773,m774,m775,m776,m777,m778,m779,m780,m781,m782,m783,n0,n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n30,n31,n32,n33,n34,n35,n36,n37,n38,n39,n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n50,n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80,n81,n82,n83,n84,n85,n86,n87,n88,n89,n90,n91,n92,n93,n94,n95,n96,n97,n98,n99,n100,n101,n102,n103,n104,n105,n106,n107,n108,n109,n110,n111,n112,n113,n114,n115,n116,n117,n118,n119,n120,n121,n122,n123,n124,n125,n126,n127,n128,n129,n130,n131,n132,n133,n134,n135,n136,n137,n138,n139,n140,n141,n142,n143,n144,n145,n146,n147,n148,n149,n150,n151,n152,n153,n154,n155,n156,n157,n158,n159,n160,n161,n162,n163,n164,n165,n166,n167,n168,n169,n170,n171,n172,n173,n174,n175,n176,n177,n178,n179,n180,n181,n182,n183,n184,n185,n186,n187,n188,n189,n190,n191,n192,n193,n194,n195,n196,n197,n198,n199,n200,n201,n202,n203,n204,n205,n206,n207,n208,n209,n210,n211,n212,n213,n214,n215,n216,n217,n218,n219,n220,n221,n222,n223,n224,n225,n226,n227,n228,n229,n230,n231,n232,n233,n234,n235,n236,n237,n238,n239,n240,n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,n251,n252,n253,n254,n255,n256,n257,n258,n259,n260,n261,n262,n263,n264,n265,n266,n267,n268,n269,n270,n271,n272,n273,n274,n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,n330,n331,n332,n333,n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,n345,n346,n347,n348,n349,n350,n351,n352,n353,n354,n355,n356,n357,n358,n359,n360,n361,n362,n363,n364,n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,n385,n386,n387,n388,n389,n390,n391,n392,n393,n394,n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,n415,n416,n417,n418,n419,n420,n421,n422,n423,n424,n425,n426,n427,n428,n429,n430,n431,n432,n433,n434,n435,n436,n437,n438,n439,n440,n441,n442,n443,n444,n445,n446,n447,n448,n449,n450,n451,n452,n453,n454,n455,n456,n457,n458,n459,n460,n461,n462,n463,n464,n465,n466,n467,n468,n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,n479,n480,n481,n482,n483,n484,n485,n486,n487,n488,n489,n490,n491,n492,n493,n494,n495,n496,n497,n498,n499,n500,n501,n502,n503,n504,n505,n506,n507,n508,n509,n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,n559,n560,n561,n562,n563,n564,n565,n566,n567,n568,n569,n570,n571,n572,n573,n574,n575,n576,n577,n578,n579,n580,n581,n582,n583,n584,n585,n586,n587,n588,n589,n590,n591,n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,n612,n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,n623,n624,n625,n626,n627,n628,n629,n630,n631,n632,n633,n634,n635,n636,n637,n638,n639,n640,n641,n642,n643,n644,n645,n646,n647,n648,n649,n650,n651,n652,n653,n654,n655,n656,n657,n658,n659,n660,n661,n662,n663,n664,n665,n666,n667,n668,n669,n670,n671,n672,n673,n674,n675,n676,n677,n678,n679,n680,n681,n682,n683,n684,n685,n686,n687,n688,n689,n690,n691,n692,n693,n694,n695,n696,n697,n698,n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,n709,n710,n711,n712,n713,n714,n715,n716,n717,n718,n719,n720,n721,n722,n723,n724,n725,n726,n727,n728,n729,n730,n731,n732,n733,n734,n735,n736,n737,n738,n739,n740,n741,n742,n743,n744,n745,n746,n747,n748,n749,n750,n751,n752,n753,n754,n755,n756,n757,n758,n759,n760,n761,n762,n763,n764,n765,n766,n767,n768,n769,n770,n771,n772,n773,n774,n775,n776,n777,n778,n779,n780,n781,n782,n783;
  
  localparam integer a0 = 0;
    generate 
        localparam integer b0 = 0;
        for (m0 = 0; m0 < 16; m0 = m0 + 1) 
        begin: inbit0
            assign data_11[m0 + b0*16 + a0*28*16] = data_11_array[a0][b0][m0];
        end
    endgenerate
    generate 
        localparam integer b1 = 1;
        for (m1 = 0; m1 < 16; m1 = m1 + 1) 
        begin: inbit1
            assign data_11[m1 + b1*16 + a0*28*16] = data_11_array[a0][b1][m1];
        end
    endgenerate
    generate 
        localparam integer b2 = 2;
        for (m2 = 0; m2 < 16; m2 = m2 + 1) 
        begin: inbit2
            assign data_11[m2 + b2*16 + a0*28*16] = data_11_array[a0][b2][m2];
        end
    endgenerate
    generate 
        localparam integer b3 = 3;
        for (m3 = 0; m3 < 16; m3 = m3 + 1) 
        begin: inbit3
            assign data_11[m3 + b3*16 + a0*28*16] = data_11_array[a0][b3][m3];
        end
    endgenerate
    generate 
        localparam integer b4 = 4;
        for (m4 = 0; m4 < 16; m4 = m4 + 1) 
        begin: inbit4
            assign data_11[m4 + b4*16 + a0*28*16] = data_11_array[a0][b4][m4];
        end
    endgenerate
    generate 
        localparam integer b5 = 5;
        for (m5 = 0; m5 < 16; m5 = m5 + 1) 
        begin: inbit5
            assign data_11[m5 + b5*16 + a0*28*16] = data_11_array[a0][b5][m5];
        end
    endgenerate
    generate 
        localparam integer b6 = 6;
        for (m6 = 0; m6 < 16; m6 = m6 + 1) 
        begin: inbit6
            assign data_11[m6 + b6*16 + a0*28*16] = data_11_array[a0][b6][m6];
        end
    endgenerate
    generate 
        localparam integer b7 = 7;
        for (m7 = 0; m7 < 16; m7 = m7 + 1) 
        begin: inbit7
            assign data_11[m7 + b7*16 + a0*28*16] = data_11_array[a0][b7][m7];
        end
    endgenerate
    generate 
        localparam integer b8 = 8;
        for (m8 = 0; m8 < 16; m8 = m8 + 1) 
        begin: inbit8
            assign data_11[m8 + b8*16 + a0*28*16] = data_11_array[a0][b8][m8];
        end
    endgenerate
    generate 
        localparam integer b9 = 9;
        for (m9 = 0; m9 < 16; m9 = m9 + 1) 
        begin: inbit9
            assign data_11[m9 + b9*16 + a0*28*16] = data_11_array[a0][b9][m9];
        end
    endgenerate
    generate 
        localparam integer b10 = 10;
        for (m10 = 0; m10 < 16; m10 = m10 + 1) 
        begin: inbit10
            assign data_11[m10 + b10*16 + a0*28*16] = data_11_array[a0][b10][m10];
        end
    endgenerate
    generate 
        localparam integer b11 = 11;
        for (m11 = 0; m11 < 16; m11 = m11 + 1) 
        begin: inbit11
            assign data_11[m11 + b11*16 + a0*28*16] = data_11_array[a0][b11][m11];
        end
    endgenerate
    generate 
        localparam integer b12 = 12;
        for (m12 = 0; m12 < 16; m12 = m12 + 1) 
        begin: inbit12
            assign data_11[m12 + b12*16 + a0*28*16] = data_11_array[a0][b12][m12];
        end
    endgenerate
    generate 
        localparam integer b13 = 13;
        for (m13 = 0; m13 < 16; m13 = m13 + 1) 
        begin: inbit13
            assign data_11[m13 + b13*16 + a0*28*16] = data_11_array[a0][b13][m13];
        end
    endgenerate
    generate 
        localparam integer b14 = 14;
        for (m14 = 0; m14 < 16; m14 = m14 + 1) 
        begin: inbit14
            assign data_11[m14 + b14*16 + a0*28*16] = data_11_array[a0][b14][m14];
        end
    endgenerate
    generate 
        localparam integer b15 = 15;
        for (m15 = 0; m15 < 16; m15 = m15 + 1) 
        begin: inbit15
            assign data_11[m15 + b15*16 + a0*28*16] = data_11_array[a0][b15][m15];
        end
    endgenerate
    generate 
        localparam integer b16 = 16;
        for (m16 = 0; m16 < 16; m16 = m16 + 1) 
        begin: inbit16
            assign data_11[m16 + b16*16 + a0*28*16] = data_11_array[a0][b16][m16];
        end
    endgenerate
    generate 
        localparam integer b17 = 17;
        for (m17 = 0; m17 < 16; m17 = m17 + 1) 
        begin: inbit17
            assign data_11[m17 + b17*16 + a0*28*16] = data_11_array[a0][b17][m17];
        end
    endgenerate
    generate 
        localparam integer b18 = 18;
        for (m18 = 0; m18 < 16; m18 = m18 + 1) 
        begin: inbit18
            assign data_11[m18 + b18*16 + a0*28*16] = data_11_array[a0][b18][m18];
        end
    endgenerate
    generate 
        localparam integer b19 = 19;
        for (m19 = 0; m19 < 16; m19 = m19 + 1) 
        begin: inbit19
            assign data_11[m19 + b19*16 + a0*28*16] = data_11_array[a0][b19][m19];
        end
    endgenerate
    generate 
        localparam integer b20 = 20;
        for (m20 = 0; m20 < 16; m20 = m20 + 1) 
        begin: inbit20
            assign data_11[m20 + b20*16 + a0*28*16] = data_11_array[a0][b20][m20];
        end
    endgenerate
    generate 
        localparam integer b21 = 21;
        for (m21 = 0; m21 < 16; m21 = m21 + 1) 
        begin: inbit21
            assign data_11[m21 + b21*16 + a0*28*16] = data_11_array[a0][b21][m21];
        end
    endgenerate
    generate 
        localparam integer b22 = 22;
        for (m22 = 0; m22 < 16; m22 = m22 + 1) 
        begin: inbit22
            assign data_11[m22 + b22*16 + a0*28*16] = data_11_array[a0][b22][m22];
        end
    endgenerate
    generate 
        localparam integer b23 = 23;
        for (m23 = 0; m23 < 16; m23 = m23 + 1) 
        begin: inbit23
            assign data_11[m23 + b23*16 + a0*28*16] = data_11_array[a0][b23][m23];
        end
    endgenerate
    generate 
        localparam integer b24 = 24;
        for (m24 = 0; m24 < 16; m24 = m24 + 1) 
        begin: inbit24
            assign data_11[m24 + b24*16 + a0*28*16] = data_11_array[a0][b24][m24];
        end
    endgenerate
    generate 
        localparam integer b25 = 25;
        for (m25 = 0; m25 < 16; m25 = m25 + 1) 
        begin: inbit25
            assign data_11[m25 + b25*16 + a0*28*16] = data_11_array[a0][b25][m25];
        end
    endgenerate
    generate 
        localparam integer b26 = 26;
        for (m26 = 0; m26 < 16; m26 = m26 + 1) 
        begin: inbit26
            assign data_11[m26 + b26*16 + a0*28*16] = data_11_array[a0][b26][m26];
        end
    endgenerate
    generate 
        localparam integer b27 = 27;
        for (m27 = 0; m27 < 16; m27 = m27 + 1) 
        begin: inbit27
            assign data_11[m27 + b27*16 + a0*28*16] = data_11_array[a0][b27][m27];
        end
    endgenerate
    localparam integer a1 = 1;
    generate 
        localparam integer b28 = 0;
        for (m28 = 0; m28 < 16; m28 = m28 + 1) 
        begin: inbit28
            assign data_11[m28 + b28*16 + a1*28*16] = data_11_array[a1][b28][m28];
        end
    endgenerate
    generate 
        localparam integer b29 = 1;
        for (m29 = 0; m29 < 16; m29 = m29 + 1) 
        begin: inbit29
            assign data_11[m29 + b29*16 + a1*28*16] = data_11_array[a1][b29][m29];
        end
    endgenerate
    generate 
        localparam integer b30 = 2;
        for (m30 = 0; m30 < 16; m30 = m30 + 1) 
        begin: inbit30
            assign data_11[m30 + b30*16 + a1*28*16] = data_11_array[a1][b30][m30];
        end
    endgenerate
    generate 
        localparam integer b31 = 3;
        for (m31 = 0; m31 < 16; m31 = m31 + 1) 
        begin: inbit31
            assign data_11[m31 + b31*16 + a1*28*16] = data_11_array[a1][b31][m31];
        end
    endgenerate
    generate 
        localparam integer b32 = 4;
        for (m32 = 0; m32 < 16; m32 = m32 + 1) 
        begin: inbit32
            assign data_11[m32 + b32*16 + a1*28*16] = data_11_array[a1][b32][m32];
        end
    endgenerate
    generate 
        localparam integer b33 = 5;
        for (m33 = 0; m33 < 16; m33 = m33 + 1) 
        begin: inbit33
            assign data_11[m33 + b33*16 + a1*28*16] = data_11_array[a1][b33][m33];
        end
    endgenerate
    generate 
        localparam integer b34 = 6;
        for (m34 = 0; m34 < 16; m34 = m34 + 1) 
        begin: inbit34
            assign data_11[m34 + b34*16 + a1*28*16] = data_11_array[a1][b34][m34];
        end
    endgenerate
    generate 
        localparam integer b35 = 7;
        for (m35 = 0; m35 < 16; m35 = m35 + 1) 
        begin: inbit35
            assign data_11[m35 + b35*16 + a1*28*16] = data_11_array[a1][b35][m35];
        end
    endgenerate
    generate 
        localparam integer b36 = 8;
        for (m36 = 0; m36 < 16; m36 = m36 + 1) 
        begin: inbit36
            assign data_11[m36 + b36*16 + a1*28*16] = data_11_array[a1][b36][m36];
        end
    endgenerate
    generate 
        localparam integer b37 = 9;
        for (m37 = 0; m37 < 16; m37 = m37 + 1) 
        begin: inbit37
            assign data_11[m37 + b37*16 + a1*28*16] = data_11_array[a1][b37][m37];
        end
    endgenerate
    generate 
        localparam integer b38 = 10;
        for (m38 = 0; m38 < 16; m38 = m38 + 1) 
        begin: inbit38
            assign data_11[m38 + b38*16 + a1*28*16] = data_11_array[a1][b38][m38];
        end
    endgenerate
    generate 
        localparam integer b39 = 11;
        for (m39 = 0; m39 < 16; m39 = m39 + 1) 
        begin: inbit39
            assign data_11[m39 + b39*16 + a1*28*16] = data_11_array[a1][b39][m39];
        end
    endgenerate
    generate 
        localparam integer b40 = 12;
        for (m40 = 0; m40 < 16; m40 = m40 + 1) 
        begin: inbit40
            assign data_11[m40 + b40*16 + a1*28*16] = data_11_array[a1][b40][m40];
        end
    endgenerate
    generate 
        localparam integer b41 = 13;
        for (m41 = 0; m41 < 16; m41 = m41 + 1) 
        begin: inbit41
            assign data_11[m41 + b41*16 + a1*28*16] = data_11_array[a1][b41][m41];
        end
    endgenerate
    generate 
        localparam integer b42 = 14;
        for (m42 = 0; m42 < 16; m42 = m42 + 1) 
        begin: inbit42
            assign data_11[m42 + b42*16 + a1*28*16] = data_11_array[a1][b42][m42];
        end
    endgenerate
    generate 
        localparam integer b43 = 15;
        for (m43 = 0; m43 < 16; m43 = m43 + 1) 
        begin: inbit43
            assign data_11[m43 + b43*16 + a1*28*16] = data_11_array[a1][b43][m43];
        end
    endgenerate
    generate 
        localparam integer b44 = 16;
        for (m44 = 0; m44 < 16; m44 = m44 + 1) 
        begin: inbit44
            assign data_11[m44 + b44*16 + a1*28*16] = data_11_array[a1][b44][m44];
        end
    endgenerate
    generate 
        localparam integer b45 = 17;
        for (m45 = 0; m45 < 16; m45 = m45 + 1) 
        begin: inbit45
            assign data_11[m45 + b45*16 + a1*28*16] = data_11_array[a1][b45][m45];
        end
    endgenerate
    generate 
        localparam integer b46 = 18;
        for (m46 = 0; m46 < 16; m46 = m46 + 1) 
        begin: inbit46
            assign data_11[m46 + b46*16 + a1*28*16] = data_11_array[a1][b46][m46];
        end
    endgenerate
    generate 
        localparam integer b47 = 19;
        for (m47 = 0; m47 < 16; m47 = m47 + 1) 
        begin: inbit47
            assign data_11[m47 + b47*16 + a1*28*16] = data_11_array[a1][b47][m47];
        end
    endgenerate
    generate 
        localparam integer b48 = 20;
        for (m48 = 0; m48 < 16; m48 = m48 + 1) 
        begin: inbit48
            assign data_11[m48 + b48*16 + a1*28*16] = data_11_array[a1][b48][m48];
        end
    endgenerate
    generate 
        localparam integer b49 = 21;
        for (m49 = 0; m49 < 16; m49 = m49 + 1) 
        begin: inbit49
            assign data_11[m49 + b49*16 + a1*28*16] = data_11_array[a1][b49][m49];
        end
    endgenerate
    generate 
        localparam integer b50 = 22;
        for (m50 = 0; m50 < 16; m50 = m50 + 1) 
        begin: inbit50
            assign data_11[m50 + b50*16 + a1*28*16] = data_11_array[a1][b50][m50];
        end
    endgenerate
    generate 
        localparam integer b51 = 23;
        for (m51 = 0; m51 < 16; m51 = m51 + 1) 
        begin: inbit51
            assign data_11[m51 + b51*16 + a1*28*16] = data_11_array[a1][b51][m51];
        end
    endgenerate
    generate 
        localparam integer b52 = 24;
        for (m52 = 0; m52 < 16; m52 = m52 + 1) 
        begin: inbit52
            assign data_11[m52 + b52*16 + a1*28*16] = data_11_array[a1][b52][m52];
        end
    endgenerate
    generate 
        localparam integer b53 = 25;
        for (m53 = 0; m53 < 16; m53 = m53 + 1) 
        begin: inbit53
            assign data_11[m53 + b53*16 + a1*28*16] = data_11_array[a1][b53][m53];
        end
    endgenerate
    generate 
        localparam integer b54 = 26;
        for (m54 = 0; m54 < 16; m54 = m54 + 1) 
        begin: inbit54
            assign data_11[m54 + b54*16 + a1*28*16] = data_11_array[a1][b54][m54];
        end
    endgenerate
    generate 
        localparam integer b55 = 27;
        for (m55 = 0; m55 < 16; m55 = m55 + 1) 
        begin: inbit55
            assign data_11[m55 + b55*16 + a1*28*16] = data_11_array[a1][b55][m55];
        end
    endgenerate
    localparam integer a2 = 2;
    generate 
        localparam integer b56 = 0;
        for (m56 = 0; m56 < 16; m56 = m56 + 1) 
        begin: inbit56
            assign data_11[m56 + b56*16 + a2*28*16] = data_11_array[a2][b56][m56];
        end
    endgenerate
    generate 
        localparam integer b57 = 1;
        for (m57 = 0; m57 < 16; m57 = m57 + 1) 
        begin: inbit57
            assign data_11[m57 + b57*16 + a2*28*16] = data_11_array[a2][b57][m57];
        end
    endgenerate
    generate 
        localparam integer b58 = 2;
        for (m58 = 0; m58 < 16; m58 = m58 + 1) 
        begin: inbit58
            assign data_11[m58 + b58*16 + a2*28*16] = data_11_array[a2][b58][m58];
        end
    endgenerate
    generate 
        localparam integer b59 = 3;
        for (m59 = 0; m59 < 16; m59 = m59 + 1) 
        begin: inbit59
            assign data_11[m59 + b59*16 + a2*28*16] = data_11_array[a2][b59][m59];
        end
    endgenerate
    generate 
        localparam integer b60 = 4;
        for (m60 = 0; m60 < 16; m60 = m60 + 1) 
        begin: inbit60
            assign data_11[m60 + b60*16 + a2*28*16] = data_11_array[a2][b60][m60];
        end
    endgenerate
    generate 
        localparam integer b61 = 5;
        for (m61 = 0; m61 < 16; m61 = m61 + 1) 
        begin: inbit61
            assign data_11[m61 + b61*16 + a2*28*16] = data_11_array[a2][b61][m61];
        end
    endgenerate
    generate 
        localparam integer b62 = 6;
        for (m62 = 0; m62 < 16; m62 = m62 + 1) 
        begin: inbit62
            assign data_11[m62 + b62*16 + a2*28*16] = data_11_array[a2][b62][m62];
        end
    endgenerate
    generate 
        localparam integer b63 = 7;
        for (m63 = 0; m63 < 16; m63 = m63 + 1) 
        begin: inbit63
            assign data_11[m63 + b63*16 + a2*28*16] = data_11_array[a2][b63][m63];
        end
    endgenerate
    generate 
        localparam integer b64 = 8;
        for (m64 = 0; m64 < 16; m64 = m64 + 1) 
        begin: inbit64
            assign data_11[m64 + b64*16 + a2*28*16] = data_11_array[a2][b64][m64];
        end
    endgenerate
    generate 
        localparam integer b65 = 9;
        for (m65 = 0; m65 < 16; m65 = m65 + 1) 
        begin: inbit65
            assign data_11[m65 + b65*16 + a2*28*16] = data_11_array[a2][b65][m65];
        end
    endgenerate
    generate 
        localparam integer b66 = 10;
        for (m66 = 0; m66 < 16; m66 = m66 + 1) 
        begin: inbit66
            assign data_11[m66 + b66*16 + a2*28*16] = data_11_array[a2][b66][m66];
        end
    endgenerate
    generate 
        localparam integer b67 = 11;
        for (m67 = 0; m67 < 16; m67 = m67 + 1) 
        begin: inbit67
            assign data_11[m67 + b67*16 + a2*28*16] = data_11_array[a2][b67][m67];
        end
    endgenerate
    generate 
        localparam integer b68 = 12;
        for (m68 = 0; m68 < 16; m68 = m68 + 1) 
        begin: inbit68
            assign data_11[m68 + b68*16 + a2*28*16] = data_11_array[a2][b68][m68];
        end
    endgenerate
    generate 
        localparam integer b69 = 13;
        for (m69 = 0; m69 < 16; m69 = m69 + 1) 
        begin: inbit69
            assign data_11[m69 + b69*16 + a2*28*16] = data_11_array[a2][b69][m69];
        end
    endgenerate
    generate 
        localparam integer b70 = 14;
        for (m70 = 0; m70 < 16; m70 = m70 + 1) 
        begin: inbit70
            assign data_11[m70 + b70*16 + a2*28*16] = data_11_array[a2][b70][m70];
        end
    endgenerate
    generate 
        localparam integer b71 = 15;
        for (m71 = 0; m71 < 16; m71 = m71 + 1) 
        begin: inbit71
            assign data_11[m71 + b71*16 + a2*28*16] = data_11_array[a2][b71][m71];
        end
    endgenerate
    generate 
        localparam integer b72 = 16;
        for (m72 = 0; m72 < 16; m72 = m72 + 1) 
        begin: inbit72
            assign data_11[m72 + b72*16 + a2*28*16] = data_11_array[a2][b72][m72];
        end
    endgenerate
    generate 
        localparam integer b73 = 17;
        for (m73 = 0; m73 < 16; m73 = m73 + 1) 
        begin: inbit73
            assign data_11[m73 + b73*16 + a2*28*16] = data_11_array[a2][b73][m73];
        end
    endgenerate
    generate 
        localparam integer b74 = 18;
        for (m74 = 0; m74 < 16; m74 = m74 + 1) 
        begin: inbit74
            assign data_11[m74 + b74*16 + a2*28*16] = data_11_array[a2][b74][m74];
        end
    endgenerate
    generate 
        localparam integer b75 = 19;
        for (m75 = 0; m75 < 16; m75 = m75 + 1) 
        begin: inbit75
            assign data_11[m75 + b75*16 + a2*28*16] = data_11_array[a2][b75][m75];
        end
    endgenerate
    generate 
        localparam integer b76 = 20;
        for (m76 = 0; m76 < 16; m76 = m76 + 1) 
        begin: inbit76
            assign data_11[m76 + b76*16 + a2*28*16] = data_11_array[a2][b76][m76];
        end
    endgenerate
    generate 
        localparam integer b77 = 21;
        for (m77 = 0; m77 < 16; m77 = m77 + 1) 
        begin: inbit77
            assign data_11[m77 + b77*16 + a2*28*16] = data_11_array[a2][b77][m77];
        end
    endgenerate
    generate 
        localparam integer b78 = 22;
        for (m78 = 0; m78 < 16; m78 = m78 + 1) 
        begin: inbit78
            assign data_11[m78 + b78*16 + a2*28*16] = data_11_array[a2][b78][m78];
        end
    endgenerate
    generate 
        localparam integer b79 = 23;
        for (m79 = 0; m79 < 16; m79 = m79 + 1) 
        begin: inbit79
            assign data_11[m79 + b79*16 + a2*28*16] = data_11_array[a2][b79][m79];
        end
    endgenerate
    generate 
        localparam integer b80 = 24;
        for (m80 = 0; m80 < 16; m80 = m80 + 1) 
        begin: inbit80
            assign data_11[m80 + b80*16 + a2*28*16] = data_11_array[a2][b80][m80];
        end
    endgenerate
    generate 
        localparam integer b81 = 25;
        for (m81 = 0; m81 < 16; m81 = m81 + 1) 
        begin: inbit81
            assign data_11[m81 + b81*16 + a2*28*16] = data_11_array[a2][b81][m81];
        end
    endgenerate
    generate 
        localparam integer b82 = 26;
        for (m82 = 0; m82 < 16; m82 = m82 + 1) 
        begin: inbit82
            assign data_11[m82 + b82*16 + a2*28*16] = data_11_array[a2][b82][m82];
        end
    endgenerate
    generate 
        localparam integer b83 = 27;
        for (m83 = 0; m83 < 16; m83 = m83 + 1) 
        begin: inbit83
            assign data_11[m83 + b83*16 + a2*28*16] = data_11_array[a2][b83][m83];
        end
    endgenerate
    localparam integer a3 = 3;
    generate 
        localparam integer b84 = 0;
        for (m84 = 0; m84 < 16; m84 = m84 + 1) 
        begin: inbit84
            assign data_11[m84 + b84*16 + a3*28*16] = data_11_array[a3][b84][m84];
        end
    endgenerate
    generate 
        localparam integer b85 = 1;
        for (m85 = 0; m85 < 16; m85 = m85 + 1) 
        begin: inbit85
            assign data_11[m85 + b85*16 + a3*28*16] = data_11_array[a3][b85][m85];
        end
    endgenerate
    generate 
        localparam integer b86 = 2;
        for (m86 = 0; m86 < 16; m86 = m86 + 1) 
        begin: inbit86
            assign data_11[m86 + b86*16 + a3*28*16] = data_11_array[a3][b86][m86];
        end
    endgenerate
    generate 
        localparam integer b87 = 3;
        for (m87 = 0; m87 < 16; m87 = m87 + 1) 
        begin: inbit87
            assign data_11[m87 + b87*16 + a3*28*16] = data_11_array[a3][b87][m87];
        end
    endgenerate
    generate 
        localparam integer b88 = 4;
        for (m88 = 0; m88 < 16; m88 = m88 + 1) 
        begin: inbit88
            assign data_11[m88 + b88*16 + a3*28*16] = data_11_array[a3][b88][m88];
        end
    endgenerate
    generate 
        localparam integer b89 = 5;
        for (m89 = 0; m89 < 16; m89 = m89 + 1) 
        begin: inbit89
            assign data_11[m89 + b89*16 + a3*28*16] = data_11_array[a3][b89][m89];
        end
    endgenerate
    generate 
        localparam integer b90 = 6;
        for (m90 = 0; m90 < 16; m90 = m90 + 1) 
        begin: inbit90
            assign data_11[m90 + b90*16 + a3*28*16] = data_11_array[a3][b90][m90];
        end
    endgenerate
    generate 
        localparam integer b91 = 7;
        for (m91 = 0; m91 < 16; m91 = m91 + 1) 
        begin: inbit91
            assign data_11[m91 + b91*16 + a3*28*16] = data_11_array[a3][b91][m91];
        end
    endgenerate
    generate 
        localparam integer b92 = 8;
        for (m92 = 0; m92 < 16; m92 = m92 + 1) 
        begin: inbit92
            assign data_11[m92 + b92*16 + a3*28*16] = data_11_array[a3][b92][m92];
        end
    endgenerate
    generate 
        localparam integer b93 = 9;
        for (m93 = 0; m93 < 16; m93 = m93 + 1) 
        begin: inbit93
            assign data_11[m93 + b93*16 + a3*28*16] = data_11_array[a3][b93][m93];
        end
    endgenerate
    generate 
        localparam integer b94 = 10;
        for (m94 = 0; m94 < 16; m94 = m94 + 1) 
        begin: inbit94
            assign data_11[m94 + b94*16 + a3*28*16] = data_11_array[a3][b94][m94];
        end
    endgenerate
    generate 
        localparam integer b95 = 11;
        for (m95 = 0; m95 < 16; m95 = m95 + 1) 
        begin: inbit95
            assign data_11[m95 + b95*16 + a3*28*16] = data_11_array[a3][b95][m95];
        end
    endgenerate
    generate 
        localparam integer b96 = 12;
        for (m96 = 0; m96 < 16; m96 = m96 + 1) 
        begin: inbit96
            assign data_11[m96 + b96*16 + a3*28*16] = data_11_array[a3][b96][m96];
        end
    endgenerate
    generate 
        localparam integer b97 = 13;
        for (m97 = 0; m97 < 16; m97 = m97 + 1) 
        begin: inbit97
            assign data_11[m97 + b97*16 + a3*28*16] = data_11_array[a3][b97][m97];
        end
    endgenerate
    generate 
        localparam integer b98 = 14;
        for (m98 = 0; m98 < 16; m98 = m98 + 1) 
        begin: inbit98
            assign data_11[m98 + b98*16 + a3*28*16] = data_11_array[a3][b98][m98];
        end
    endgenerate
    generate 
        localparam integer b99 = 15;
        for (m99 = 0; m99 < 16; m99 = m99 + 1) 
        begin: inbit99
            assign data_11[m99 + b99*16 + a3*28*16] = data_11_array[a3][b99][m99];
        end
    endgenerate
    generate 
        localparam integer b100 = 16;
        for (m100 = 0; m100 < 16; m100 = m100 + 1) 
        begin: inbit100
            assign data_11[m100 + b100*16 + a3*28*16] = data_11_array[a3][b100][m100];
        end
    endgenerate
    generate 
        localparam integer b101 = 17;
        for (m101 = 0; m101 < 16; m101 = m101 + 1) 
        begin: inbit101
            assign data_11[m101 + b101*16 + a3*28*16] = data_11_array[a3][b101][m101];
        end
    endgenerate
    generate 
        localparam integer b102 = 18;
        for (m102 = 0; m102 < 16; m102 = m102 + 1) 
        begin: inbit102
            assign data_11[m102 + b102*16 + a3*28*16] = data_11_array[a3][b102][m102];
        end
    endgenerate
    generate 
        localparam integer b103 = 19;
        for (m103 = 0; m103 < 16; m103 = m103 + 1) 
        begin: inbit103
            assign data_11[m103 + b103*16 + a3*28*16] = data_11_array[a3][b103][m103];
        end
    endgenerate
    generate 
        localparam integer b104 = 20;
        for (m104 = 0; m104 < 16; m104 = m104 + 1) 
        begin: inbit104
            assign data_11[m104 + b104*16 + a3*28*16] = data_11_array[a3][b104][m104];
        end
    endgenerate
    generate 
        localparam integer b105 = 21;
        for (m105 = 0; m105 < 16; m105 = m105 + 1) 
        begin: inbit105
            assign data_11[m105 + b105*16 + a3*28*16] = data_11_array[a3][b105][m105];
        end
    endgenerate
    generate 
        localparam integer b106 = 22;
        for (m106 = 0; m106 < 16; m106 = m106 + 1) 
        begin: inbit106
            assign data_11[m106 + b106*16 + a3*28*16] = data_11_array[a3][b106][m106];
        end
    endgenerate
    generate 
        localparam integer b107 = 23;
        for (m107 = 0; m107 < 16; m107 = m107 + 1) 
        begin: inbit107
            assign data_11[m107 + b107*16 + a3*28*16] = data_11_array[a3][b107][m107];
        end
    endgenerate
    generate 
        localparam integer b108 = 24;
        for (m108 = 0; m108 < 16; m108 = m108 + 1) 
        begin: inbit108
            assign data_11[m108 + b108*16 + a3*28*16] = data_11_array[a3][b108][m108];
        end
    endgenerate
    generate 
        localparam integer b109 = 25;
        for (m109 = 0; m109 < 16; m109 = m109 + 1) 
        begin: inbit109
            assign data_11[m109 + b109*16 + a3*28*16] = data_11_array[a3][b109][m109];
        end
    endgenerate
    generate 
        localparam integer b110 = 26;
        for (m110 = 0; m110 < 16; m110 = m110 + 1) 
        begin: inbit110
            assign data_11[m110 + b110*16 + a3*28*16] = data_11_array[a3][b110][m110];
        end
    endgenerate
    generate 
        localparam integer b111 = 27;
        for (m111 = 0; m111 < 16; m111 = m111 + 1) 
        begin: inbit111
            assign data_11[m111 + b111*16 + a3*28*16] = data_11_array[a3][b111][m111];
        end
    endgenerate
    localparam integer a4 = 4;
    generate 
        localparam integer b112 = 0;
        for (m112 = 0; m112 < 16; m112 = m112 + 1) 
        begin: inbit112
            assign data_11[m112 + b112*16 + a4*28*16] = data_11_array[a4][b112][m112];
        end
    endgenerate
    generate 
        localparam integer b113 = 1;
        for (m113 = 0; m113 < 16; m113 = m113 + 1) 
        begin: inbit113
            assign data_11[m113 + b113*16 + a4*28*16] = data_11_array[a4][b113][m113];
        end
    endgenerate
    generate 
        localparam integer b114 = 2;
        for (m114 = 0; m114 < 16; m114 = m114 + 1) 
        begin: inbit114
            assign data_11[m114 + b114*16 + a4*28*16] = data_11_array[a4][b114][m114];
        end
    endgenerate
    generate 
        localparam integer b115 = 3;
        for (m115 = 0; m115 < 16; m115 = m115 + 1) 
        begin: inbit115
            assign data_11[m115 + b115*16 + a4*28*16] = data_11_array[a4][b115][m115];
        end
    endgenerate
    generate 
        localparam integer b116 = 4;
        for (m116 = 0; m116 < 16; m116 = m116 + 1) 
        begin: inbit116
            assign data_11[m116 + b116*16 + a4*28*16] = data_11_array[a4][b116][m116];
        end
    endgenerate
    generate 
        localparam integer b117 = 5;
        for (m117 = 0; m117 < 16; m117 = m117 + 1) 
        begin: inbit117
            assign data_11[m117 + b117*16 + a4*28*16] = data_11_array[a4][b117][m117];
        end
    endgenerate
    generate 
        localparam integer b118 = 6;
        for (m118 = 0; m118 < 16; m118 = m118 + 1) 
        begin: inbit118
            assign data_11[m118 + b118*16 + a4*28*16] = data_11_array[a4][b118][m118];
        end
    endgenerate
    generate 
        localparam integer b119 = 7;
        for (m119 = 0; m119 < 16; m119 = m119 + 1) 
        begin: inbit119
            assign data_11[m119 + b119*16 + a4*28*16] = data_11_array[a4][b119][m119];
        end
    endgenerate
    generate 
        localparam integer b120 = 8;
        for (m120 = 0; m120 < 16; m120 = m120 + 1) 
        begin: inbit120
            assign data_11[m120 + b120*16 + a4*28*16] = data_11_array[a4][b120][m120];
        end
    endgenerate
    generate 
        localparam integer b121 = 9;
        for (m121 = 0; m121 < 16; m121 = m121 + 1) 
        begin: inbit121
            assign data_11[m121 + b121*16 + a4*28*16] = data_11_array[a4][b121][m121];
        end
    endgenerate
    generate 
        localparam integer b122 = 10;
        for (m122 = 0; m122 < 16; m122 = m122 + 1) 
        begin: inbit122
            assign data_11[m122 + b122*16 + a4*28*16] = data_11_array[a4][b122][m122];
        end
    endgenerate
    generate 
        localparam integer b123 = 11;
        for (m123 = 0; m123 < 16; m123 = m123 + 1) 
        begin: inbit123
            assign data_11[m123 + b123*16 + a4*28*16] = data_11_array[a4][b123][m123];
        end
    endgenerate
    generate 
        localparam integer b124 = 12;
        for (m124 = 0; m124 < 16; m124 = m124 + 1) 
        begin: inbit124
            assign data_11[m124 + b124*16 + a4*28*16] = data_11_array[a4][b124][m124];
        end
    endgenerate
    generate 
        localparam integer b125 = 13;
        for (m125 = 0; m125 < 16; m125 = m125 + 1) 
        begin: inbit125
            assign data_11[m125 + b125*16 + a4*28*16] = data_11_array[a4][b125][m125];
        end
    endgenerate
    generate 
        localparam integer b126 = 14;
        for (m126 = 0; m126 < 16; m126 = m126 + 1) 
        begin: inbit126
            assign data_11[m126 + b126*16 + a4*28*16] = data_11_array[a4][b126][m126];
        end
    endgenerate
    generate 
        localparam integer b127 = 15;
        for (m127 = 0; m127 < 16; m127 = m127 + 1) 
        begin: inbit127
            assign data_11[m127 + b127*16 + a4*28*16] = data_11_array[a4][b127][m127];
        end
    endgenerate
    generate 
        localparam integer b128 = 16;
        for (m128 = 0; m128 < 16; m128 = m128 + 1) 
        begin: inbit128
            assign data_11[m128 + b128*16 + a4*28*16] = data_11_array[a4][b128][m128];
        end
    endgenerate
    generate 
        localparam integer b129 = 17;
        for (m129 = 0; m129 < 16; m129 = m129 + 1) 
        begin: inbit129
            assign data_11[m129 + b129*16 + a4*28*16] = data_11_array[a4][b129][m129];
        end
    endgenerate
    generate 
        localparam integer b130 = 18;
        for (m130 = 0; m130 < 16; m130 = m130 + 1) 
        begin: inbit130
            assign data_11[m130 + b130*16 + a4*28*16] = data_11_array[a4][b130][m130];
        end
    endgenerate
    generate 
        localparam integer b131 = 19;
        for (m131 = 0; m131 < 16; m131 = m131 + 1) 
        begin: inbit131
            assign data_11[m131 + b131*16 + a4*28*16] = data_11_array[a4][b131][m131];
        end
    endgenerate
    generate 
        localparam integer b132 = 20;
        for (m132 = 0; m132 < 16; m132 = m132 + 1) 
        begin: inbit132
            assign data_11[m132 + b132*16 + a4*28*16] = data_11_array[a4][b132][m132];
        end
    endgenerate
    generate 
        localparam integer b133 = 21;
        for (m133 = 0; m133 < 16; m133 = m133 + 1) 
        begin: inbit133
            assign data_11[m133 + b133*16 + a4*28*16] = data_11_array[a4][b133][m133];
        end
    endgenerate
    generate 
        localparam integer b134 = 22;
        for (m134 = 0; m134 < 16; m134 = m134 + 1) 
        begin: inbit134
            assign data_11[m134 + b134*16 + a4*28*16] = data_11_array[a4][b134][m134];
        end
    endgenerate
    generate 
        localparam integer b135 = 23;
        for (m135 = 0; m135 < 16; m135 = m135 + 1) 
        begin: inbit135
            assign data_11[m135 + b135*16 + a4*28*16] = data_11_array[a4][b135][m135];
        end
    endgenerate
    generate 
        localparam integer b136 = 24;
        for (m136 = 0; m136 < 16; m136 = m136 + 1) 
        begin: inbit136
            assign data_11[m136 + b136*16 + a4*28*16] = data_11_array[a4][b136][m136];
        end
    endgenerate
    generate 
        localparam integer b137 = 25;
        for (m137 = 0; m137 < 16; m137 = m137 + 1) 
        begin: inbit137
            assign data_11[m137 + b137*16 + a4*28*16] = data_11_array[a4][b137][m137];
        end
    endgenerate
    generate 
        localparam integer b138 = 26;
        for (m138 = 0; m138 < 16; m138 = m138 + 1) 
        begin: inbit138
            assign data_11[m138 + b138*16 + a4*28*16] = data_11_array[a4][b138][m138];
        end
    endgenerate
    generate 
        localparam integer b139 = 27;
        for (m139 = 0; m139 < 16; m139 = m139 + 1) 
        begin: inbit139
            assign data_11[m139 + b139*16 + a4*28*16] = data_11_array[a4][b139][m139];
        end
    endgenerate
    localparam integer a5 = 5;
    generate 
        localparam integer b140 = 0;
        for (m140 = 0; m140 < 16; m140 = m140 + 1) 
        begin: inbit140
            assign data_11[m140 + b140*16 + a5*28*16] = data_11_array[a5][b140][m140];
        end
    endgenerate
    generate 
        localparam integer b141 = 1;
        for (m141 = 0; m141 < 16; m141 = m141 + 1) 
        begin: inbit141
            assign data_11[m141 + b141*16 + a5*28*16] = data_11_array[a5][b141][m141];
        end
    endgenerate
    generate 
        localparam integer b142 = 2;
        for (m142 = 0; m142 < 16; m142 = m142 + 1) 
        begin: inbit142
            assign data_11[m142 + b142*16 + a5*28*16] = data_11_array[a5][b142][m142];
        end
    endgenerate
    generate 
        localparam integer b143 = 3;
        for (m143 = 0; m143 < 16; m143 = m143 + 1) 
        begin: inbit143
            assign data_11[m143 + b143*16 + a5*28*16] = data_11_array[a5][b143][m143];
        end
    endgenerate
    generate 
        localparam integer b144 = 4;
        for (m144 = 0; m144 < 16; m144 = m144 + 1) 
        begin: inbit144
            assign data_11[m144 + b144*16 + a5*28*16] = data_11_array[a5][b144][m144];
        end
    endgenerate
    generate 
        localparam integer b145 = 5;
        for (m145 = 0; m145 < 16; m145 = m145 + 1) 
        begin: inbit145
            assign data_11[m145 + b145*16 + a5*28*16] = data_11_array[a5][b145][m145];
        end
    endgenerate
    generate 
        localparam integer b146 = 6;
        for (m146 = 0; m146 < 16; m146 = m146 + 1) 
        begin: inbit146
            assign data_11[m146 + b146*16 + a5*28*16] = data_11_array[a5][b146][m146];
        end
    endgenerate
    generate 
        localparam integer b147 = 7;
        for (m147 = 0; m147 < 16; m147 = m147 + 1) 
        begin: inbit147
            assign data_11[m147 + b147*16 + a5*28*16] = data_11_array[a5][b147][m147];
        end
    endgenerate
    generate 
        localparam integer b148 = 8;
        for (m148 = 0; m148 < 16; m148 = m148 + 1) 
        begin: inbit148
            assign data_11[m148 + b148*16 + a5*28*16] = data_11_array[a5][b148][m148];
        end
    endgenerate
    generate 
        localparam integer b149 = 9;
        for (m149 = 0; m149 < 16; m149 = m149 + 1) 
        begin: inbit149
            assign data_11[m149 + b149*16 + a5*28*16] = data_11_array[a5][b149][m149];
        end
    endgenerate
    generate 
        localparam integer b150 = 10;
        for (m150 = 0; m150 < 16; m150 = m150 + 1) 
        begin: inbit150
            assign data_11[m150 + b150*16 + a5*28*16] = data_11_array[a5][b150][m150];
        end
    endgenerate
    generate 
        localparam integer b151 = 11;
        for (m151 = 0; m151 < 16; m151 = m151 + 1) 
        begin: inbit151
            assign data_11[m151 + b151*16 + a5*28*16] = data_11_array[a5][b151][m151];
        end
    endgenerate
    generate 
        localparam integer b152 = 12;
        for (m152 = 0; m152 < 16; m152 = m152 + 1) 
        begin: inbit152
            assign data_11[m152 + b152*16 + a5*28*16] = data_11_array[a5][b152][m152];
        end
    endgenerate
    generate 
        localparam integer b153 = 13;
        for (m153 = 0; m153 < 16; m153 = m153 + 1) 
        begin: inbit153
            assign data_11[m153 + b153*16 + a5*28*16] = data_11_array[a5][b153][m153];
        end
    endgenerate
    generate 
        localparam integer b154 = 14;
        for (m154 = 0; m154 < 16; m154 = m154 + 1) 
        begin: inbit154
            assign data_11[m154 + b154*16 + a5*28*16] = data_11_array[a5][b154][m154];
        end
    endgenerate
    generate 
        localparam integer b155 = 15;
        for (m155 = 0; m155 < 16; m155 = m155 + 1) 
        begin: inbit155
            assign data_11[m155 + b155*16 + a5*28*16] = data_11_array[a5][b155][m155];
        end
    endgenerate
    generate 
        localparam integer b156 = 16;
        for (m156 = 0; m156 < 16; m156 = m156 + 1) 
        begin: inbit156
            assign data_11[m156 + b156*16 + a5*28*16] = data_11_array[a5][b156][m156];
        end
    endgenerate
    generate 
        localparam integer b157 = 17;
        for (m157 = 0; m157 < 16; m157 = m157 + 1) 
        begin: inbit157
            assign data_11[m157 + b157*16 + a5*28*16] = data_11_array[a5][b157][m157];
        end
    endgenerate
    generate 
        localparam integer b158 = 18;
        for (m158 = 0; m158 < 16; m158 = m158 + 1) 
        begin: inbit158
            assign data_11[m158 + b158*16 + a5*28*16] = data_11_array[a5][b158][m158];
        end
    endgenerate
    generate 
        localparam integer b159 = 19;
        for (m159 = 0; m159 < 16; m159 = m159 + 1) 
        begin: inbit159
            assign data_11[m159 + b159*16 + a5*28*16] = data_11_array[a5][b159][m159];
        end
    endgenerate
    generate 
        localparam integer b160 = 20;
        for (m160 = 0; m160 < 16; m160 = m160 + 1) 
        begin: inbit160
            assign data_11[m160 + b160*16 + a5*28*16] = data_11_array[a5][b160][m160];
        end
    endgenerate
    generate 
        localparam integer b161 = 21;
        for (m161 = 0; m161 < 16; m161 = m161 + 1) 
        begin: inbit161
            assign data_11[m161 + b161*16 + a5*28*16] = data_11_array[a5][b161][m161];
        end
    endgenerate
    generate 
        localparam integer b162 = 22;
        for (m162 = 0; m162 < 16; m162 = m162 + 1) 
        begin: inbit162
            assign data_11[m162 + b162*16 + a5*28*16] = data_11_array[a5][b162][m162];
        end
    endgenerate
    generate 
        localparam integer b163 = 23;
        for (m163 = 0; m163 < 16; m163 = m163 + 1) 
        begin: inbit163
            assign data_11[m163 + b163*16 + a5*28*16] = data_11_array[a5][b163][m163];
        end
    endgenerate
    generate 
        localparam integer b164 = 24;
        for (m164 = 0; m164 < 16; m164 = m164 + 1) 
        begin: inbit164
            assign data_11[m164 + b164*16 + a5*28*16] = data_11_array[a5][b164][m164];
        end
    endgenerate
    generate 
        localparam integer b165 = 25;
        for (m165 = 0; m165 < 16; m165 = m165 + 1) 
        begin: inbit165
            assign data_11[m165 + b165*16 + a5*28*16] = data_11_array[a5][b165][m165];
        end
    endgenerate
    generate 
        localparam integer b166 = 26;
        for (m166 = 0; m166 < 16; m166 = m166 + 1) 
        begin: inbit166
            assign data_11[m166 + b166*16 + a5*28*16] = data_11_array[a5][b166][m166];
        end
    endgenerate
    generate 
        localparam integer b167 = 27;
        for (m167 = 0; m167 < 16; m167 = m167 + 1) 
        begin: inbit167
            assign data_11[m167 + b167*16 + a5*28*16] = data_11_array[a5][b167][m167];
        end
    endgenerate
    localparam integer a6 = 6;
    generate 
        localparam integer b168 = 0;
        for (m168 = 0; m168 < 16; m168 = m168 + 1) 
        begin: inbit168
            assign data_11[m168 + b168*16 + a6*28*16] = data_11_array[a6][b168][m168];
        end
    endgenerate
    generate 
        localparam integer b169 = 1;
        for (m169 = 0; m169 < 16; m169 = m169 + 1) 
        begin: inbit169
            assign data_11[m169 + b169*16 + a6*28*16] = data_11_array[a6][b169][m169];
        end
    endgenerate
    generate 
        localparam integer b170 = 2;
        for (m170 = 0; m170 < 16; m170 = m170 + 1) 
        begin: inbit170
            assign data_11[m170 + b170*16 + a6*28*16] = data_11_array[a6][b170][m170];
        end
    endgenerate
    generate 
        localparam integer b171 = 3;
        for (m171 = 0; m171 < 16; m171 = m171 + 1) 
        begin: inbit171
            assign data_11[m171 + b171*16 + a6*28*16] = data_11_array[a6][b171][m171];
        end
    endgenerate
    generate 
        localparam integer b172 = 4;
        for (m172 = 0; m172 < 16; m172 = m172 + 1) 
        begin: inbit172
            assign data_11[m172 + b172*16 + a6*28*16] = data_11_array[a6][b172][m172];
        end
    endgenerate
    generate 
        localparam integer b173 = 5;
        for (m173 = 0; m173 < 16; m173 = m173 + 1) 
        begin: inbit173
            assign data_11[m173 + b173*16 + a6*28*16] = data_11_array[a6][b173][m173];
        end
    endgenerate
    generate 
        localparam integer b174 = 6;
        for (m174 = 0; m174 < 16; m174 = m174 + 1) 
        begin: inbit174
            assign data_11[m174 + b174*16 + a6*28*16] = data_11_array[a6][b174][m174];
        end
    endgenerate
    generate 
        localparam integer b175 = 7;
        for (m175 = 0; m175 < 16; m175 = m175 + 1) 
        begin: inbit175
            assign data_11[m175 + b175*16 + a6*28*16] = data_11_array[a6][b175][m175];
        end
    endgenerate
    generate 
        localparam integer b176 = 8;
        for (m176 = 0; m176 < 16; m176 = m176 + 1) 
        begin: inbit176
            assign data_11[m176 + b176*16 + a6*28*16] = data_11_array[a6][b176][m176];
        end
    endgenerate
    generate 
        localparam integer b177 = 9;
        for (m177 = 0; m177 < 16; m177 = m177 + 1) 
        begin: inbit177
            assign data_11[m177 + b177*16 + a6*28*16] = data_11_array[a6][b177][m177];
        end
    endgenerate
    generate 
        localparam integer b178 = 10;
        for (m178 = 0; m178 < 16; m178 = m178 + 1) 
        begin: inbit178
            assign data_11[m178 + b178*16 + a6*28*16] = data_11_array[a6][b178][m178];
        end
    endgenerate
    generate 
        localparam integer b179 = 11;
        for (m179 = 0; m179 < 16; m179 = m179 + 1) 
        begin: inbit179
            assign data_11[m179 + b179*16 + a6*28*16] = data_11_array[a6][b179][m179];
        end
    endgenerate
    generate 
        localparam integer b180 = 12;
        for (m180 = 0; m180 < 16; m180 = m180 + 1) 
        begin: inbit180
            assign data_11[m180 + b180*16 + a6*28*16] = data_11_array[a6][b180][m180];
        end
    endgenerate
    generate 
        localparam integer b181 = 13;
        for (m181 = 0; m181 < 16; m181 = m181 + 1) 
        begin: inbit181
            assign data_11[m181 + b181*16 + a6*28*16] = data_11_array[a6][b181][m181];
        end
    endgenerate
    generate 
        localparam integer b182 = 14;
        for (m182 = 0; m182 < 16; m182 = m182 + 1) 
        begin: inbit182
            assign data_11[m182 + b182*16 + a6*28*16] = data_11_array[a6][b182][m182];
        end
    endgenerate
    generate 
        localparam integer b183 = 15;
        for (m183 = 0; m183 < 16; m183 = m183 + 1) 
        begin: inbit183
            assign data_11[m183 + b183*16 + a6*28*16] = data_11_array[a6][b183][m183];
        end
    endgenerate
    generate 
        localparam integer b184 = 16;
        for (m184 = 0; m184 < 16; m184 = m184 + 1) 
        begin: inbit184
            assign data_11[m184 + b184*16 + a6*28*16] = data_11_array[a6][b184][m184];
        end
    endgenerate
    generate 
        localparam integer b185 = 17;
        for (m185 = 0; m185 < 16; m185 = m185 + 1) 
        begin: inbit185
            assign data_11[m185 + b185*16 + a6*28*16] = data_11_array[a6][b185][m185];
        end
    endgenerate
    generate 
        localparam integer b186 = 18;
        for (m186 = 0; m186 < 16; m186 = m186 + 1) 
        begin: inbit186
            assign data_11[m186 + b186*16 + a6*28*16] = data_11_array[a6][b186][m186];
        end
    endgenerate
    generate 
        localparam integer b187 = 19;
        for (m187 = 0; m187 < 16; m187 = m187 + 1) 
        begin: inbit187
            assign data_11[m187 + b187*16 + a6*28*16] = data_11_array[a6][b187][m187];
        end
    endgenerate
    generate 
        localparam integer b188 = 20;
        for (m188 = 0; m188 < 16; m188 = m188 + 1) 
        begin: inbit188
            assign data_11[m188 + b188*16 + a6*28*16] = data_11_array[a6][b188][m188];
        end
    endgenerate
    generate 
        localparam integer b189 = 21;
        for (m189 = 0; m189 < 16; m189 = m189 + 1) 
        begin: inbit189
            assign data_11[m189 + b189*16 + a6*28*16] = data_11_array[a6][b189][m189];
        end
    endgenerate
    generate 
        localparam integer b190 = 22;
        for (m190 = 0; m190 < 16; m190 = m190 + 1) 
        begin: inbit190
            assign data_11[m190 + b190*16 + a6*28*16] = data_11_array[a6][b190][m190];
        end
    endgenerate
    generate 
        localparam integer b191 = 23;
        for (m191 = 0; m191 < 16; m191 = m191 + 1) 
        begin: inbit191
            assign data_11[m191 + b191*16 + a6*28*16] = data_11_array[a6][b191][m191];
        end
    endgenerate
    generate 
        localparam integer b192 = 24;
        for (m192 = 0; m192 < 16; m192 = m192 + 1) 
        begin: inbit192
            assign data_11[m192 + b192*16 + a6*28*16] = data_11_array[a6][b192][m192];
        end
    endgenerate
    generate 
        localparam integer b193 = 25;
        for (m193 = 0; m193 < 16; m193 = m193 + 1) 
        begin: inbit193
            assign data_11[m193 + b193*16 + a6*28*16] = data_11_array[a6][b193][m193];
        end
    endgenerate
    generate 
        localparam integer b194 = 26;
        for (m194 = 0; m194 < 16; m194 = m194 + 1) 
        begin: inbit194
            assign data_11[m194 + b194*16 + a6*28*16] = data_11_array[a6][b194][m194];
        end
    endgenerate
    generate 
        localparam integer b195 = 27;
        for (m195 = 0; m195 < 16; m195 = m195 + 1) 
        begin: inbit195
            assign data_11[m195 + b195*16 + a6*28*16] = data_11_array[a6][b195][m195];
        end
    endgenerate
    localparam integer a7 = 7;
    generate 
        localparam integer b196 = 0;
        for (m196 = 0; m196 < 16; m196 = m196 + 1) 
        begin: inbit196
            assign data_11[m196 + b196*16 + a7*28*16] = data_11_array[a7][b196][m196];
        end
    endgenerate
    generate 
        localparam integer b197 = 1;
        for (m197 = 0; m197 < 16; m197 = m197 + 1) 
        begin: inbit197
            assign data_11[m197 + b197*16 + a7*28*16] = data_11_array[a7][b197][m197];
        end
    endgenerate
    generate 
        localparam integer b198 = 2;
        for (m198 = 0; m198 < 16; m198 = m198 + 1) 
        begin: inbit198
            assign data_11[m198 + b198*16 + a7*28*16] = data_11_array[a7][b198][m198];
        end
    endgenerate
    generate 
        localparam integer b199 = 3;
        for (m199 = 0; m199 < 16; m199 = m199 + 1) 
        begin: inbit199
            assign data_11[m199 + b199*16 + a7*28*16] = data_11_array[a7][b199][m199];
        end
    endgenerate
    generate 
        localparam integer b200 = 4;
        for (m200 = 0; m200 < 16; m200 = m200 + 1) 
        begin: inbit200
            assign data_11[m200 + b200*16 + a7*28*16] = data_11_array[a7][b200][m200];
        end
    endgenerate
    generate 
        localparam integer b201 = 5;
        for (m201 = 0; m201 < 16; m201 = m201 + 1) 
        begin: inbit201
            assign data_11[m201 + b201*16 + a7*28*16] = data_11_array[a7][b201][m201];
        end
    endgenerate
    generate 
        localparam integer b202 = 6;
        for (m202 = 0; m202 < 16; m202 = m202 + 1) 
        begin: inbit202
            assign data_11[m202 + b202*16 + a7*28*16] = data_11_array[a7][b202][m202];
        end
    endgenerate
    generate 
        localparam integer b203 = 7;
        for (m203 = 0; m203 < 16; m203 = m203 + 1) 
        begin: inbit203
            assign data_11[m203 + b203*16 + a7*28*16] = data_11_array[a7][b203][m203];
        end
    endgenerate
    generate 
        localparam integer b204 = 8;
        for (m204 = 0; m204 < 16; m204 = m204 + 1) 
        begin: inbit204
            assign data_11[m204 + b204*16 + a7*28*16] = data_11_array[a7][b204][m204];
        end
    endgenerate
    generate 
        localparam integer b205 = 9;
        for (m205 = 0; m205 < 16; m205 = m205 + 1) 
        begin: inbit205
            assign data_11[m205 + b205*16 + a7*28*16] = data_11_array[a7][b205][m205];
        end
    endgenerate
    generate 
        localparam integer b206 = 10;
        for (m206 = 0; m206 < 16; m206 = m206 + 1) 
        begin: inbit206
            assign data_11[m206 + b206*16 + a7*28*16] = data_11_array[a7][b206][m206];
        end
    endgenerate
    generate 
        localparam integer b207 = 11;
        for (m207 = 0; m207 < 16; m207 = m207 + 1) 
        begin: inbit207
            assign data_11[m207 + b207*16 + a7*28*16] = data_11_array[a7][b207][m207];
        end
    endgenerate
    generate 
        localparam integer b208 = 12;
        for (m208 = 0; m208 < 16; m208 = m208 + 1) 
        begin: inbit208
            assign data_11[m208 + b208*16 + a7*28*16] = data_11_array[a7][b208][m208];
        end
    endgenerate
    generate 
        localparam integer b209 = 13;
        for (m209 = 0; m209 < 16; m209 = m209 + 1) 
        begin: inbit209
            assign data_11[m209 + b209*16 + a7*28*16] = data_11_array[a7][b209][m209];
        end
    endgenerate
    generate 
        localparam integer b210 = 14;
        for (m210 = 0; m210 < 16; m210 = m210 + 1) 
        begin: inbit210
            assign data_11[m210 + b210*16 + a7*28*16] = data_11_array[a7][b210][m210];
        end
    endgenerate
    generate 
        localparam integer b211 = 15;
        for (m211 = 0; m211 < 16; m211 = m211 + 1) 
        begin: inbit211
            assign data_11[m211 + b211*16 + a7*28*16] = data_11_array[a7][b211][m211];
        end
    endgenerate
    generate 
        localparam integer b212 = 16;
        for (m212 = 0; m212 < 16; m212 = m212 + 1) 
        begin: inbit212
            assign data_11[m212 + b212*16 + a7*28*16] = data_11_array[a7][b212][m212];
        end
    endgenerate
    generate 
        localparam integer b213 = 17;
        for (m213 = 0; m213 < 16; m213 = m213 + 1) 
        begin: inbit213
            assign data_11[m213 + b213*16 + a7*28*16] = data_11_array[a7][b213][m213];
        end
    endgenerate
    generate 
        localparam integer b214 = 18;
        for (m214 = 0; m214 < 16; m214 = m214 + 1) 
        begin: inbit214
            assign data_11[m214 + b214*16 + a7*28*16] = data_11_array[a7][b214][m214];
        end
    endgenerate
    generate 
        localparam integer b215 = 19;
        for (m215 = 0; m215 < 16; m215 = m215 + 1) 
        begin: inbit215
            assign data_11[m215 + b215*16 + a7*28*16] = data_11_array[a7][b215][m215];
        end
    endgenerate
    generate 
        localparam integer b216 = 20;
        for (m216 = 0; m216 < 16; m216 = m216 + 1) 
        begin: inbit216
            assign data_11[m216 + b216*16 + a7*28*16] = data_11_array[a7][b216][m216];
        end
    endgenerate
    generate 
        localparam integer b217 = 21;
        for (m217 = 0; m217 < 16; m217 = m217 + 1) 
        begin: inbit217
            assign data_11[m217 + b217*16 + a7*28*16] = data_11_array[a7][b217][m217];
        end
    endgenerate
    generate 
        localparam integer b218 = 22;
        for (m218 = 0; m218 < 16; m218 = m218 + 1) 
        begin: inbit218
            assign data_11[m218 + b218*16 + a7*28*16] = data_11_array[a7][b218][m218];
        end
    endgenerate
    generate 
        localparam integer b219 = 23;
        for (m219 = 0; m219 < 16; m219 = m219 + 1) 
        begin: inbit219
            assign data_11[m219 + b219*16 + a7*28*16] = data_11_array[a7][b219][m219];
        end
    endgenerate
    generate 
        localparam integer b220 = 24;
        for (m220 = 0; m220 < 16; m220 = m220 + 1) 
        begin: inbit220
            assign data_11[m220 + b220*16 + a7*28*16] = data_11_array[a7][b220][m220];
        end
    endgenerate
    generate 
        localparam integer b221 = 25;
        for (m221 = 0; m221 < 16; m221 = m221 + 1) 
        begin: inbit221
            assign data_11[m221 + b221*16 + a7*28*16] = data_11_array[a7][b221][m221];
        end
    endgenerate
    generate 
        localparam integer b222 = 26;
        for (m222 = 0; m222 < 16; m222 = m222 + 1) 
        begin: inbit222
            assign data_11[m222 + b222*16 + a7*28*16] = data_11_array[a7][b222][m222];
        end
    endgenerate
    generate 
        localparam integer b223 = 27;
        for (m223 = 0; m223 < 16; m223 = m223 + 1) 
        begin: inbit223
            assign data_11[m223 + b223*16 + a7*28*16] = data_11_array[a7][b223][m223];
        end
    endgenerate
    localparam integer a8 = 8;
    generate 
        localparam integer b224 = 0;
        for (m224 = 0; m224 < 16; m224 = m224 + 1) 
        begin: inbit224
            assign data_11[m224 + b224*16 + a8*28*16] = data_11_array[a8][b224][m224];
        end
    endgenerate
    generate 
        localparam integer b225 = 1;
        for (m225 = 0; m225 < 16; m225 = m225 + 1) 
        begin: inbit225
            assign data_11[m225 + b225*16 + a8*28*16] = data_11_array[a8][b225][m225];
        end
    endgenerate
    generate 
        localparam integer b226 = 2;
        for (m226 = 0; m226 < 16; m226 = m226 + 1) 
        begin: inbit226
            assign data_11[m226 + b226*16 + a8*28*16] = data_11_array[a8][b226][m226];
        end
    endgenerate
    generate 
        localparam integer b227 = 3;
        for (m227 = 0; m227 < 16; m227 = m227 + 1) 
        begin: inbit227
            assign data_11[m227 + b227*16 + a8*28*16] = data_11_array[a8][b227][m227];
        end
    endgenerate
    generate 
        localparam integer b228 = 4;
        for (m228 = 0; m228 < 16; m228 = m228 + 1) 
        begin: inbit228
            assign data_11[m228 + b228*16 + a8*28*16] = data_11_array[a8][b228][m228];
        end
    endgenerate
    generate 
        localparam integer b229 = 5;
        for (m229 = 0; m229 < 16; m229 = m229 + 1) 
        begin: inbit229
            assign data_11[m229 + b229*16 + a8*28*16] = data_11_array[a8][b229][m229];
        end
    endgenerate
    generate 
        localparam integer b230 = 6;
        for (m230 = 0; m230 < 16; m230 = m230 + 1) 
        begin: inbit230
            assign data_11[m230 + b230*16 + a8*28*16] = data_11_array[a8][b230][m230];
        end
    endgenerate
    generate 
        localparam integer b231 = 7;
        for (m231 = 0; m231 < 16; m231 = m231 + 1) 
        begin: inbit231
            assign data_11[m231 + b231*16 + a8*28*16] = data_11_array[a8][b231][m231];
        end
    endgenerate
    generate 
        localparam integer b232 = 8;
        for (m232 = 0; m232 < 16; m232 = m232 + 1) 
        begin: inbit232
            assign data_11[m232 + b232*16 + a8*28*16] = data_11_array[a8][b232][m232];
        end
    endgenerate
    generate 
        localparam integer b233 = 9;
        for (m233 = 0; m233 < 16; m233 = m233 + 1) 
        begin: inbit233
            assign data_11[m233 + b233*16 + a8*28*16] = data_11_array[a8][b233][m233];
        end
    endgenerate
    generate 
        localparam integer b234 = 10;
        for (m234 = 0; m234 < 16; m234 = m234 + 1) 
        begin: inbit234
            assign data_11[m234 + b234*16 + a8*28*16] = data_11_array[a8][b234][m234];
        end
    endgenerate
    generate 
        localparam integer b235 = 11;
        for (m235 = 0; m235 < 16; m235 = m235 + 1) 
        begin: inbit235
            assign data_11[m235 + b235*16 + a8*28*16] = data_11_array[a8][b235][m235];
        end
    endgenerate
    generate 
        localparam integer b236 = 12;
        for (m236 = 0; m236 < 16; m236 = m236 + 1) 
        begin: inbit236
            assign data_11[m236 + b236*16 + a8*28*16] = data_11_array[a8][b236][m236];
        end
    endgenerate
    generate 
        localparam integer b237 = 13;
        for (m237 = 0; m237 < 16; m237 = m237 + 1) 
        begin: inbit237
            assign data_11[m237 + b237*16 + a8*28*16] = data_11_array[a8][b237][m237];
        end
    endgenerate
    generate 
        localparam integer b238 = 14;
        for (m238 = 0; m238 < 16; m238 = m238 + 1) 
        begin: inbit238
            assign data_11[m238 + b238*16 + a8*28*16] = data_11_array[a8][b238][m238];
        end
    endgenerate
    generate 
        localparam integer b239 = 15;
        for (m239 = 0; m239 < 16; m239 = m239 + 1) 
        begin: inbit239
            assign data_11[m239 + b239*16 + a8*28*16] = data_11_array[a8][b239][m239];
        end
    endgenerate
    generate 
        localparam integer b240 = 16;
        for (m240 = 0; m240 < 16; m240 = m240 + 1) 
        begin: inbit240
            assign data_11[m240 + b240*16 + a8*28*16] = data_11_array[a8][b240][m240];
        end
    endgenerate
    generate 
        localparam integer b241 = 17;
        for (m241 = 0; m241 < 16; m241 = m241 + 1) 
        begin: inbit241
            assign data_11[m241 + b241*16 + a8*28*16] = data_11_array[a8][b241][m241];
        end
    endgenerate
    generate 
        localparam integer b242 = 18;
        for (m242 = 0; m242 < 16; m242 = m242 + 1) 
        begin: inbit242
            assign data_11[m242 + b242*16 + a8*28*16] = data_11_array[a8][b242][m242];
        end
    endgenerate
    generate 
        localparam integer b243 = 19;
        for (m243 = 0; m243 < 16; m243 = m243 + 1) 
        begin: inbit243
            assign data_11[m243 + b243*16 + a8*28*16] = data_11_array[a8][b243][m243];
        end
    endgenerate
    generate 
        localparam integer b244 = 20;
        for (m244 = 0; m244 < 16; m244 = m244 + 1) 
        begin: inbit244
            assign data_11[m244 + b244*16 + a8*28*16] = data_11_array[a8][b244][m244];
        end
    endgenerate
    generate 
        localparam integer b245 = 21;
        for (m245 = 0; m245 < 16; m245 = m245 + 1) 
        begin: inbit245
            assign data_11[m245 + b245*16 + a8*28*16] = data_11_array[a8][b245][m245];
        end
    endgenerate
    generate 
        localparam integer b246 = 22;
        for (m246 = 0; m246 < 16; m246 = m246 + 1) 
        begin: inbit246
            assign data_11[m246 + b246*16 + a8*28*16] = data_11_array[a8][b246][m246];
        end
    endgenerate
    generate 
        localparam integer b247 = 23;
        for (m247 = 0; m247 < 16; m247 = m247 + 1) 
        begin: inbit247
            assign data_11[m247 + b247*16 + a8*28*16] = data_11_array[a8][b247][m247];
        end
    endgenerate
    generate 
        localparam integer b248 = 24;
        for (m248 = 0; m248 < 16; m248 = m248 + 1) 
        begin: inbit248
            assign data_11[m248 + b248*16 + a8*28*16] = data_11_array[a8][b248][m248];
        end
    endgenerate
    generate 
        localparam integer b249 = 25;
        for (m249 = 0; m249 < 16; m249 = m249 + 1) 
        begin: inbit249
            assign data_11[m249 + b249*16 + a8*28*16] = data_11_array[a8][b249][m249];
        end
    endgenerate
    generate 
        localparam integer b250 = 26;
        for (m250 = 0; m250 < 16; m250 = m250 + 1) 
        begin: inbit250
            assign data_11[m250 + b250*16 + a8*28*16] = data_11_array[a8][b250][m250];
        end
    endgenerate
    generate 
        localparam integer b251 = 27;
        for (m251 = 0; m251 < 16; m251 = m251 + 1) 
        begin: inbit251
            assign data_11[m251 + b251*16 + a8*28*16] = data_11_array[a8][b251][m251];
        end
    endgenerate
    localparam integer a9 = 9;
    generate 
        localparam integer b252 = 0;
        for (m252 = 0; m252 < 16; m252 = m252 + 1) 
        begin: inbit252
            assign data_11[m252 + b252*16 + a9*28*16] = data_11_array[a9][b252][m252];
        end
    endgenerate
    generate 
        localparam integer b253 = 1;
        for (m253 = 0; m253 < 16; m253 = m253 + 1) 
        begin: inbit253
            assign data_11[m253 + b253*16 + a9*28*16] = data_11_array[a9][b253][m253];
        end
    endgenerate
    generate 
        localparam integer b254 = 2;
        for (m254 = 0; m254 < 16; m254 = m254 + 1) 
        begin: inbit254
            assign data_11[m254 + b254*16 + a9*28*16] = data_11_array[a9][b254][m254];
        end
    endgenerate
    generate 
        localparam integer b255 = 3;
        for (m255 = 0; m255 < 16; m255 = m255 + 1) 
        begin: inbit255
            assign data_11[m255 + b255*16 + a9*28*16] = data_11_array[a9][b255][m255];
        end
    endgenerate
    generate 
        localparam integer b256 = 4;
        for (m256 = 0; m256 < 16; m256 = m256 + 1) 
        begin: inbit256
            assign data_11[m256 + b256*16 + a9*28*16] = data_11_array[a9][b256][m256];
        end
    endgenerate
    generate 
        localparam integer b257 = 5;
        for (m257 = 0; m257 < 16; m257 = m257 + 1) 
        begin: inbit257
            assign data_11[m257 + b257*16 + a9*28*16] = data_11_array[a9][b257][m257];
        end
    endgenerate
    generate 
        localparam integer b258 = 6;
        for (m258 = 0; m258 < 16; m258 = m258 + 1) 
        begin: inbit258
            assign data_11[m258 + b258*16 + a9*28*16] = data_11_array[a9][b258][m258];
        end
    endgenerate
    generate 
        localparam integer b259 = 7;
        for (m259 = 0; m259 < 16; m259 = m259 + 1) 
        begin: inbit259
            assign data_11[m259 + b259*16 + a9*28*16] = data_11_array[a9][b259][m259];
        end
    endgenerate
    generate 
        localparam integer b260 = 8;
        for (m260 = 0; m260 < 16; m260 = m260 + 1) 
        begin: inbit260
            assign data_11[m260 + b260*16 + a9*28*16] = data_11_array[a9][b260][m260];
        end
    endgenerate
    generate 
        localparam integer b261 = 9;
        for (m261 = 0; m261 < 16; m261 = m261 + 1) 
        begin: inbit261
            assign data_11[m261 + b261*16 + a9*28*16] = data_11_array[a9][b261][m261];
        end
    endgenerate
    generate 
        localparam integer b262 = 10;
        for (m262 = 0; m262 < 16; m262 = m262 + 1) 
        begin: inbit262
            assign data_11[m262 + b262*16 + a9*28*16] = data_11_array[a9][b262][m262];
        end
    endgenerate
    generate 
        localparam integer b263 = 11;
        for (m263 = 0; m263 < 16; m263 = m263 + 1) 
        begin: inbit263
            assign data_11[m263 + b263*16 + a9*28*16] = data_11_array[a9][b263][m263];
        end
    endgenerate
    generate 
        localparam integer b264 = 12;
        for (m264 = 0; m264 < 16; m264 = m264 + 1) 
        begin: inbit264
            assign data_11[m264 + b264*16 + a9*28*16] = data_11_array[a9][b264][m264];
        end
    endgenerate
    generate 
        localparam integer b265 = 13;
        for (m265 = 0; m265 < 16; m265 = m265 + 1) 
        begin: inbit265
            assign data_11[m265 + b265*16 + a9*28*16] = data_11_array[a9][b265][m265];
        end
    endgenerate
    generate 
        localparam integer b266 = 14;
        for (m266 = 0; m266 < 16; m266 = m266 + 1) 
        begin: inbit266
            assign data_11[m266 + b266*16 + a9*28*16] = data_11_array[a9][b266][m266];
        end
    endgenerate
    generate 
        localparam integer b267 = 15;
        for (m267 = 0; m267 < 16; m267 = m267 + 1) 
        begin: inbit267
            assign data_11[m267 + b267*16 + a9*28*16] = data_11_array[a9][b267][m267];
        end
    endgenerate
    generate 
        localparam integer b268 = 16;
        for (m268 = 0; m268 < 16; m268 = m268 + 1) 
        begin: inbit268
            assign data_11[m268 + b268*16 + a9*28*16] = data_11_array[a9][b268][m268];
        end
    endgenerate
    generate 
        localparam integer b269 = 17;
        for (m269 = 0; m269 < 16; m269 = m269 + 1) 
        begin: inbit269
            assign data_11[m269 + b269*16 + a9*28*16] = data_11_array[a9][b269][m269];
        end
    endgenerate
    generate 
        localparam integer b270 = 18;
        for (m270 = 0; m270 < 16; m270 = m270 + 1) 
        begin: inbit270
            assign data_11[m270 + b270*16 + a9*28*16] = data_11_array[a9][b270][m270];
        end
    endgenerate
    generate 
        localparam integer b271 = 19;
        for (m271 = 0; m271 < 16; m271 = m271 + 1) 
        begin: inbit271
            assign data_11[m271 + b271*16 + a9*28*16] = data_11_array[a9][b271][m271];
        end
    endgenerate
    generate 
        localparam integer b272 = 20;
        for (m272 = 0; m272 < 16; m272 = m272 + 1) 
        begin: inbit272
            assign data_11[m272 + b272*16 + a9*28*16] = data_11_array[a9][b272][m272];
        end
    endgenerate
    generate 
        localparam integer b273 = 21;
        for (m273 = 0; m273 < 16; m273 = m273 + 1) 
        begin: inbit273
            assign data_11[m273 + b273*16 + a9*28*16] = data_11_array[a9][b273][m273];
        end
    endgenerate
    generate 
        localparam integer b274 = 22;
        for (m274 = 0; m274 < 16; m274 = m274 + 1) 
        begin: inbit274
            assign data_11[m274 + b274*16 + a9*28*16] = data_11_array[a9][b274][m274];
        end
    endgenerate
    generate 
        localparam integer b275 = 23;
        for (m275 = 0; m275 < 16; m275 = m275 + 1) 
        begin: inbit275
            assign data_11[m275 + b275*16 + a9*28*16] = data_11_array[a9][b275][m275];
        end
    endgenerate
    generate 
        localparam integer b276 = 24;
        for (m276 = 0; m276 < 16; m276 = m276 + 1) 
        begin: inbit276
            assign data_11[m276 + b276*16 + a9*28*16] = data_11_array[a9][b276][m276];
        end
    endgenerate
    generate 
        localparam integer b277 = 25;
        for (m277 = 0; m277 < 16; m277 = m277 + 1) 
        begin: inbit277
            assign data_11[m277 + b277*16 + a9*28*16] = data_11_array[a9][b277][m277];
        end
    endgenerate
    generate 
        localparam integer b278 = 26;
        for (m278 = 0; m278 < 16; m278 = m278 + 1) 
        begin: inbit278
            assign data_11[m278 + b278*16 + a9*28*16] = data_11_array[a9][b278][m278];
        end
    endgenerate
    generate 
        localparam integer b279 = 27;
        for (m279 = 0; m279 < 16; m279 = m279 + 1) 
        begin: inbit279
            assign data_11[m279 + b279*16 + a9*28*16] = data_11_array[a9][b279][m279];
        end
    endgenerate
    localparam integer a10 = 10;
    generate 
        localparam integer b280 = 0;
        for (m280 = 0; m280 < 16; m280 = m280 + 1) 
        begin: inbit280
            assign data_11[m280 + b280*16 + a10*28*16] = data_11_array[a10][b280][m280];
        end
    endgenerate
    generate 
        localparam integer b281 = 1;
        for (m281 = 0; m281 < 16; m281 = m281 + 1) 
        begin: inbit281
            assign data_11[m281 + b281*16 + a10*28*16] = data_11_array[a10][b281][m281];
        end
    endgenerate
    generate 
        localparam integer b282 = 2;
        for (m282 = 0; m282 < 16; m282 = m282 + 1) 
        begin: inbit282
            assign data_11[m282 + b282*16 + a10*28*16] = data_11_array[a10][b282][m282];
        end
    endgenerate
    generate 
        localparam integer b283 = 3;
        for (m283 = 0; m283 < 16; m283 = m283 + 1) 
        begin: inbit283
            assign data_11[m283 + b283*16 + a10*28*16] = data_11_array[a10][b283][m283];
        end
    endgenerate
    generate 
        localparam integer b284 = 4;
        for (m284 = 0; m284 < 16; m284 = m284 + 1) 
        begin: inbit284
            assign data_11[m284 + b284*16 + a10*28*16] = data_11_array[a10][b284][m284];
        end
    endgenerate
    generate 
        localparam integer b285 = 5;
        for (m285 = 0; m285 < 16; m285 = m285 + 1) 
        begin: inbit285
            assign data_11[m285 + b285*16 + a10*28*16] = data_11_array[a10][b285][m285];
        end
    endgenerate
    generate 
        localparam integer b286 = 6;
        for (m286 = 0; m286 < 16; m286 = m286 + 1) 
        begin: inbit286
            assign data_11[m286 + b286*16 + a10*28*16] = data_11_array[a10][b286][m286];
        end
    endgenerate
    generate 
        localparam integer b287 = 7;
        for (m287 = 0; m287 < 16; m287 = m287 + 1) 
        begin: inbit287
            assign data_11[m287 + b287*16 + a10*28*16] = data_11_array[a10][b287][m287];
        end
    endgenerate
    generate 
        localparam integer b288 = 8;
        for (m288 = 0; m288 < 16; m288 = m288 + 1) 
        begin: inbit288
            assign data_11[m288 + b288*16 + a10*28*16] = data_11_array[a10][b288][m288];
        end
    endgenerate
    generate 
        localparam integer b289 = 9;
        for (m289 = 0; m289 < 16; m289 = m289 + 1) 
        begin: inbit289
            assign data_11[m289 + b289*16 + a10*28*16] = data_11_array[a10][b289][m289];
        end
    endgenerate
    generate 
        localparam integer b290 = 10;
        for (m290 = 0; m290 < 16; m290 = m290 + 1) 
        begin: inbit290
            assign data_11[m290 + b290*16 + a10*28*16] = data_11_array[a10][b290][m290];
        end
    endgenerate
    generate 
        localparam integer b291 = 11;
        for (m291 = 0; m291 < 16; m291 = m291 + 1) 
        begin: inbit291
            assign data_11[m291 + b291*16 + a10*28*16] = data_11_array[a10][b291][m291];
        end
    endgenerate
    generate 
        localparam integer b292 = 12;
        for (m292 = 0; m292 < 16; m292 = m292 + 1) 
        begin: inbit292
            assign data_11[m292 + b292*16 + a10*28*16] = data_11_array[a10][b292][m292];
        end
    endgenerate
    generate 
        localparam integer b293 = 13;
        for (m293 = 0; m293 < 16; m293 = m293 + 1) 
        begin: inbit293
            assign data_11[m293 + b293*16 + a10*28*16] = data_11_array[a10][b293][m293];
        end
    endgenerate
    generate 
        localparam integer b294 = 14;
        for (m294 = 0; m294 < 16; m294 = m294 + 1) 
        begin: inbit294
            assign data_11[m294 + b294*16 + a10*28*16] = data_11_array[a10][b294][m294];
        end
    endgenerate
    generate 
        localparam integer b295 = 15;
        for (m295 = 0; m295 < 16; m295 = m295 + 1) 
        begin: inbit295
            assign data_11[m295 + b295*16 + a10*28*16] = data_11_array[a10][b295][m295];
        end
    endgenerate
    generate 
        localparam integer b296 = 16;
        for (m296 = 0; m296 < 16; m296 = m296 + 1) 
        begin: inbit296
            assign data_11[m296 + b296*16 + a10*28*16] = data_11_array[a10][b296][m296];
        end
    endgenerate
    generate 
        localparam integer b297 = 17;
        for (m297 = 0; m297 < 16; m297 = m297 + 1) 
        begin: inbit297
            assign data_11[m297 + b297*16 + a10*28*16] = data_11_array[a10][b297][m297];
        end
    endgenerate
    generate 
        localparam integer b298 = 18;
        for (m298 = 0; m298 < 16; m298 = m298 + 1) 
        begin: inbit298
            assign data_11[m298 + b298*16 + a10*28*16] = data_11_array[a10][b298][m298];
        end
    endgenerate
    generate 
        localparam integer b299 = 19;
        for (m299 = 0; m299 < 16; m299 = m299 + 1) 
        begin: inbit299
            assign data_11[m299 + b299*16 + a10*28*16] = data_11_array[a10][b299][m299];
        end
    endgenerate
    generate 
        localparam integer b300 = 20;
        for (m300 = 0; m300 < 16; m300 = m300 + 1) 
        begin: inbit300
            assign data_11[m300 + b300*16 + a10*28*16] = data_11_array[a10][b300][m300];
        end
    endgenerate
    generate 
        localparam integer b301 = 21;
        for (m301 = 0; m301 < 16; m301 = m301 + 1) 
        begin: inbit301
            assign data_11[m301 + b301*16 + a10*28*16] = data_11_array[a10][b301][m301];
        end
    endgenerate
    generate 
        localparam integer b302 = 22;
        for (m302 = 0; m302 < 16; m302 = m302 + 1) 
        begin: inbit302
            assign data_11[m302 + b302*16 + a10*28*16] = data_11_array[a10][b302][m302];
        end
    endgenerate
    generate 
        localparam integer b303 = 23;
        for (m303 = 0; m303 < 16; m303 = m303 + 1) 
        begin: inbit303
            assign data_11[m303 + b303*16 + a10*28*16] = data_11_array[a10][b303][m303];
        end
    endgenerate
    generate 
        localparam integer b304 = 24;
        for (m304 = 0; m304 < 16; m304 = m304 + 1) 
        begin: inbit304
            assign data_11[m304 + b304*16 + a10*28*16] = data_11_array[a10][b304][m304];
        end
    endgenerate
    generate 
        localparam integer b305 = 25;
        for (m305 = 0; m305 < 16; m305 = m305 + 1) 
        begin: inbit305
            assign data_11[m305 + b305*16 + a10*28*16] = data_11_array[a10][b305][m305];
        end
    endgenerate
    generate 
        localparam integer b306 = 26;
        for (m306 = 0; m306 < 16; m306 = m306 + 1) 
        begin: inbit306
            assign data_11[m306 + b306*16 + a10*28*16] = data_11_array[a10][b306][m306];
        end
    endgenerate
    generate 
        localparam integer b307 = 27;
        for (m307 = 0; m307 < 16; m307 = m307 + 1) 
        begin: inbit307
            assign data_11[m307 + b307*16 + a10*28*16] = data_11_array[a10][b307][m307];
        end
    endgenerate
    localparam integer a11 = 11;
    generate 
        localparam integer b308 = 0;
        for (m308 = 0; m308 < 16; m308 = m308 + 1) 
        begin: inbit308
            assign data_11[m308 + b308*16 + a11*28*16] = data_11_array[a11][b308][m308];
        end
    endgenerate
    generate 
        localparam integer b309 = 1;
        for (m309 = 0; m309 < 16; m309 = m309 + 1) 
        begin: inbit309
            assign data_11[m309 + b309*16 + a11*28*16] = data_11_array[a11][b309][m309];
        end
    endgenerate
    generate 
        localparam integer b310 = 2;
        for (m310 = 0; m310 < 16; m310 = m310 + 1) 
        begin: inbit310
            assign data_11[m310 + b310*16 + a11*28*16] = data_11_array[a11][b310][m310];
        end
    endgenerate
    generate 
        localparam integer b311 = 3;
        for (m311 = 0; m311 < 16; m311 = m311 + 1) 
        begin: inbit311
            assign data_11[m311 + b311*16 + a11*28*16] = data_11_array[a11][b311][m311];
        end
    endgenerate
    generate 
        localparam integer b312 = 4;
        for (m312 = 0; m312 < 16; m312 = m312 + 1) 
        begin: inbit312
            assign data_11[m312 + b312*16 + a11*28*16] = data_11_array[a11][b312][m312];
        end
    endgenerate
    generate 
        localparam integer b313 = 5;
        for (m313 = 0; m313 < 16; m313 = m313 + 1) 
        begin: inbit313
            assign data_11[m313 + b313*16 + a11*28*16] = data_11_array[a11][b313][m313];
        end
    endgenerate
    generate 
        localparam integer b314 = 6;
        for (m314 = 0; m314 < 16; m314 = m314 + 1) 
        begin: inbit314
            assign data_11[m314 + b314*16 + a11*28*16] = data_11_array[a11][b314][m314];
        end
    endgenerate
    generate 
        localparam integer b315 = 7;
        for (m315 = 0; m315 < 16; m315 = m315 + 1) 
        begin: inbit315
            assign data_11[m315 + b315*16 + a11*28*16] = data_11_array[a11][b315][m315];
        end
    endgenerate
    generate 
        localparam integer b316 = 8;
        for (m316 = 0; m316 < 16; m316 = m316 + 1) 
        begin: inbit316
            assign data_11[m316 + b316*16 + a11*28*16] = data_11_array[a11][b316][m316];
        end
    endgenerate
    generate 
        localparam integer b317 = 9;
        for (m317 = 0; m317 < 16; m317 = m317 + 1) 
        begin: inbit317
            assign data_11[m317 + b317*16 + a11*28*16] = data_11_array[a11][b317][m317];
        end
    endgenerate
    generate 
        localparam integer b318 = 10;
        for (m318 = 0; m318 < 16; m318 = m318 + 1) 
        begin: inbit318
            assign data_11[m318 + b318*16 + a11*28*16] = data_11_array[a11][b318][m318];
        end
    endgenerate
    generate 
        localparam integer b319 = 11;
        for (m319 = 0; m319 < 16; m319 = m319 + 1) 
        begin: inbit319
            assign data_11[m319 + b319*16 + a11*28*16] = data_11_array[a11][b319][m319];
        end
    endgenerate
    generate 
        localparam integer b320 = 12;
        for (m320 = 0; m320 < 16; m320 = m320 + 1) 
        begin: inbit320
            assign data_11[m320 + b320*16 + a11*28*16] = data_11_array[a11][b320][m320];
        end
    endgenerate
    generate 
        localparam integer b321 = 13;
        for (m321 = 0; m321 < 16; m321 = m321 + 1) 
        begin: inbit321
            assign data_11[m321 + b321*16 + a11*28*16] = data_11_array[a11][b321][m321];
        end
    endgenerate
    generate 
        localparam integer b322 = 14;
        for (m322 = 0; m322 < 16; m322 = m322 + 1) 
        begin: inbit322
            assign data_11[m322 + b322*16 + a11*28*16] = data_11_array[a11][b322][m322];
        end
    endgenerate
    generate 
        localparam integer b323 = 15;
        for (m323 = 0; m323 < 16; m323 = m323 + 1) 
        begin: inbit323
            assign data_11[m323 + b323*16 + a11*28*16] = data_11_array[a11][b323][m323];
        end
    endgenerate
    generate 
        localparam integer b324 = 16;
        for (m324 = 0; m324 < 16; m324 = m324 + 1) 
        begin: inbit324
            assign data_11[m324 + b324*16 + a11*28*16] = data_11_array[a11][b324][m324];
        end
    endgenerate
    generate 
        localparam integer b325 = 17;
        for (m325 = 0; m325 < 16; m325 = m325 + 1) 
        begin: inbit325
            assign data_11[m325 + b325*16 + a11*28*16] = data_11_array[a11][b325][m325];
        end
    endgenerate
    generate 
        localparam integer b326 = 18;
        for (m326 = 0; m326 < 16; m326 = m326 + 1) 
        begin: inbit326
            assign data_11[m326 + b326*16 + a11*28*16] = data_11_array[a11][b326][m326];
        end
    endgenerate
    generate 
        localparam integer b327 = 19;
        for (m327 = 0; m327 < 16; m327 = m327 + 1) 
        begin: inbit327
            assign data_11[m327 + b327*16 + a11*28*16] = data_11_array[a11][b327][m327];
        end
    endgenerate
    generate 
        localparam integer b328 = 20;
        for (m328 = 0; m328 < 16; m328 = m328 + 1) 
        begin: inbit328
            assign data_11[m328 + b328*16 + a11*28*16] = data_11_array[a11][b328][m328];
        end
    endgenerate
    generate 
        localparam integer b329 = 21;
        for (m329 = 0; m329 < 16; m329 = m329 + 1) 
        begin: inbit329
            assign data_11[m329 + b329*16 + a11*28*16] = data_11_array[a11][b329][m329];
        end
    endgenerate
    generate 
        localparam integer b330 = 22;
        for (m330 = 0; m330 < 16; m330 = m330 + 1) 
        begin: inbit330
            assign data_11[m330 + b330*16 + a11*28*16] = data_11_array[a11][b330][m330];
        end
    endgenerate
    generate 
        localparam integer b331 = 23;
        for (m331 = 0; m331 < 16; m331 = m331 + 1) 
        begin: inbit331
            assign data_11[m331 + b331*16 + a11*28*16] = data_11_array[a11][b331][m331];
        end
    endgenerate
    generate 
        localparam integer b332 = 24;
        for (m332 = 0; m332 < 16; m332 = m332 + 1) 
        begin: inbit332
            assign data_11[m332 + b332*16 + a11*28*16] = data_11_array[a11][b332][m332];
        end
    endgenerate
    generate 
        localparam integer b333 = 25;
        for (m333 = 0; m333 < 16; m333 = m333 + 1) 
        begin: inbit333
            assign data_11[m333 + b333*16 + a11*28*16] = data_11_array[a11][b333][m333];
        end
    endgenerate
    generate 
        localparam integer b334 = 26;
        for (m334 = 0; m334 < 16; m334 = m334 + 1) 
        begin: inbit334
            assign data_11[m334 + b334*16 + a11*28*16] = data_11_array[a11][b334][m334];
        end
    endgenerate
    generate 
        localparam integer b335 = 27;
        for (m335 = 0; m335 < 16; m335 = m335 + 1) 
        begin: inbit335
            assign data_11[m335 + b335*16 + a11*28*16] = data_11_array[a11][b335][m335];
        end
    endgenerate
    localparam integer a12 = 12;
    generate 
        localparam integer b336 = 0;
        for (m336 = 0; m336 < 16; m336 = m336 + 1) 
        begin: inbit336
            assign data_11[m336 + b336*16 + a12*28*16] = data_11_array[a12][b336][m336];
        end
    endgenerate
    generate 
        localparam integer b337 = 1;
        for (m337 = 0; m337 < 16; m337 = m337 + 1) 
        begin: inbit337
            assign data_11[m337 + b337*16 + a12*28*16] = data_11_array[a12][b337][m337];
        end
    endgenerate
    generate 
        localparam integer b338 = 2;
        for (m338 = 0; m338 < 16; m338 = m338 + 1) 
        begin: inbit338
            assign data_11[m338 + b338*16 + a12*28*16] = data_11_array[a12][b338][m338];
        end
    endgenerate
    generate 
        localparam integer b339 = 3;
        for (m339 = 0; m339 < 16; m339 = m339 + 1) 
        begin: inbit339
            assign data_11[m339 + b339*16 + a12*28*16] = data_11_array[a12][b339][m339];
        end
    endgenerate
    generate 
        localparam integer b340 = 4;
        for (m340 = 0; m340 < 16; m340 = m340 + 1) 
        begin: inbit340
            assign data_11[m340 + b340*16 + a12*28*16] = data_11_array[a12][b340][m340];
        end
    endgenerate
    generate 
        localparam integer b341 = 5;
        for (m341 = 0; m341 < 16; m341 = m341 + 1) 
        begin: inbit341
            assign data_11[m341 + b341*16 + a12*28*16] = data_11_array[a12][b341][m341];
        end
    endgenerate
    generate 
        localparam integer b342 = 6;
        for (m342 = 0; m342 < 16; m342 = m342 + 1) 
        begin: inbit342
            assign data_11[m342 + b342*16 + a12*28*16] = data_11_array[a12][b342][m342];
        end
    endgenerate
    generate 
        localparam integer b343 = 7;
        for (m343 = 0; m343 < 16; m343 = m343 + 1) 
        begin: inbit343
            assign data_11[m343 + b343*16 + a12*28*16] = data_11_array[a12][b343][m343];
        end
    endgenerate
    generate 
        localparam integer b344 = 8;
        for (m344 = 0; m344 < 16; m344 = m344 + 1) 
        begin: inbit344
            assign data_11[m344 + b344*16 + a12*28*16] = data_11_array[a12][b344][m344];
        end
    endgenerate
    generate 
        localparam integer b345 = 9;
        for (m345 = 0; m345 < 16; m345 = m345 + 1) 
        begin: inbit345
            assign data_11[m345 + b345*16 + a12*28*16] = data_11_array[a12][b345][m345];
        end
    endgenerate
    generate 
        localparam integer b346 = 10;
        for (m346 = 0; m346 < 16; m346 = m346 + 1) 
        begin: inbit346
            assign data_11[m346 + b346*16 + a12*28*16] = data_11_array[a12][b346][m346];
        end
    endgenerate
    generate 
        localparam integer b347 = 11;
        for (m347 = 0; m347 < 16; m347 = m347 + 1) 
        begin: inbit347
            assign data_11[m347 + b347*16 + a12*28*16] = data_11_array[a12][b347][m347];
        end
    endgenerate
    generate 
        localparam integer b348 = 12;
        for (m348 = 0; m348 < 16; m348 = m348 + 1) 
        begin: inbit348
            assign data_11[m348 + b348*16 + a12*28*16] = data_11_array[a12][b348][m348];
        end
    endgenerate
    generate 
        localparam integer b349 = 13;
        for (m349 = 0; m349 < 16; m349 = m349 + 1) 
        begin: inbit349
            assign data_11[m349 + b349*16 + a12*28*16] = data_11_array[a12][b349][m349];
        end
    endgenerate
    generate 
        localparam integer b350 = 14;
        for (m350 = 0; m350 < 16; m350 = m350 + 1) 
        begin: inbit350
            assign data_11[m350 + b350*16 + a12*28*16] = data_11_array[a12][b350][m350];
        end
    endgenerate
    generate 
        localparam integer b351 = 15;
        for (m351 = 0; m351 < 16; m351 = m351 + 1) 
        begin: inbit351
            assign data_11[m351 + b351*16 + a12*28*16] = data_11_array[a12][b351][m351];
        end
    endgenerate
    generate 
        localparam integer b352 = 16;
        for (m352 = 0; m352 < 16; m352 = m352 + 1) 
        begin: inbit352
            assign data_11[m352 + b352*16 + a12*28*16] = data_11_array[a12][b352][m352];
        end
    endgenerate
    generate 
        localparam integer b353 = 17;
        for (m353 = 0; m353 < 16; m353 = m353 + 1) 
        begin: inbit353
            assign data_11[m353 + b353*16 + a12*28*16] = data_11_array[a12][b353][m353];
        end
    endgenerate
    generate 
        localparam integer b354 = 18;
        for (m354 = 0; m354 < 16; m354 = m354 + 1) 
        begin: inbit354
            assign data_11[m354 + b354*16 + a12*28*16] = data_11_array[a12][b354][m354];
        end
    endgenerate
    generate 
        localparam integer b355 = 19;
        for (m355 = 0; m355 < 16; m355 = m355 + 1) 
        begin: inbit355
            assign data_11[m355 + b355*16 + a12*28*16] = data_11_array[a12][b355][m355];
        end
    endgenerate
    generate 
        localparam integer b356 = 20;
        for (m356 = 0; m356 < 16; m356 = m356 + 1) 
        begin: inbit356
            assign data_11[m356 + b356*16 + a12*28*16] = data_11_array[a12][b356][m356];
        end
    endgenerate
    generate 
        localparam integer b357 = 21;
        for (m357 = 0; m357 < 16; m357 = m357 + 1) 
        begin: inbit357
            assign data_11[m357 + b357*16 + a12*28*16] = data_11_array[a12][b357][m357];
        end
    endgenerate
    generate 
        localparam integer b358 = 22;
        for (m358 = 0; m358 < 16; m358 = m358 + 1) 
        begin: inbit358
            assign data_11[m358 + b358*16 + a12*28*16] = data_11_array[a12][b358][m358];
        end
    endgenerate
    generate 
        localparam integer b359 = 23;
        for (m359 = 0; m359 < 16; m359 = m359 + 1) 
        begin: inbit359
            assign data_11[m359 + b359*16 + a12*28*16] = data_11_array[a12][b359][m359];
        end
    endgenerate
    generate 
        localparam integer b360 = 24;
        for (m360 = 0; m360 < 16; m360 = m360 + 1) 
        begin: inbit360
            assign data_11[m360 + b360*16 + a12*28*16] = data_11_array[a12][b360][m360];
        end
    endgenerate
    generate 
        localparam integer b361 = 25;
        for (m361 = 0; m361 < 16; m361 = m361 + 1) 
        begin: inbit361
            assign data_11[m361 + b361*16 + a12*28*16] = data_11_array[a12][b361][m361];
        end
    endgenerate
    generate 
        localparam integer b362 = 26;
        for (m362 = 0; m362 < 16; m362 = m362 + 1) 
        begin: inbit362
            assign data_11[m362 + b362*16 + a12*28*16] = data_11_array[a12][b362][m362];
        end
    endgenerate
    generate 
        localparam integer b363 = 27;
        for (m363 = 0; m363 < 16; m363 = m363 + 1) 
        begin: inbit363
            assign data_11[m363 + b363*16 + a12*28*16] = data_11_array[a12][b363][m363];
        end
    endgenerate
    localparam integer a13 = 13;
    generate 
        localparam integer b364 = 0;
        for (m364 = 0; m364 < 16; m364 = m364 + 1) 
        begin: inbit364
            assign data_11[m364 + b364*16 + a13*28*16] = data_11_array[a13][b364][m364];
        end
    endgenerate
    generate 
        localparam integer b365 = 1;
        for (m365 = 0; m365 < 16; m365 = m365 + 1) 
        begin: inbit365
            assign data_11[m365 + b365*16 + a13*28*16] = data_11_array[a13][b365][m365];
        end
    endgenerate
    generate 
        localparam integer b366 = 2;
        for (m366 = 0; m366 < 16; m366 = m366 + 1) 
        begin: inbit366
            assign data_11[m366 + b366*16 + a13*28*16] = data_11_array[a13][b366][m366];
        end
    endgenerate
    generate 
        localparam integer b367 = 3;
        for (m367 = 0; m367 < 16; m367 = m367 + 1) 
        begin: inbit367
            assign data_11[m367 + b367*16 + a13*28*16] = data_11_array[a13][b367][m367];
        end
    endgenerate
    generate 
        localparam integer b368 = 4;
        for (m368 = 0; m368 < 16; m368 = m368 + 1) 
        begin: inbit368
            assign data_11[m368 + b368*16 + a13*28*16] = data_11_array[a13][b368][m368];
        end
    endgenerate
    generate 
        localparam integer b369 = 5;
        for (m369 = 0; m369 < 16; m369 = m369 + 1) 
        begin: inbit369
            assign data_11[m369 + b369*16 + a13*28*16] = data_11_array[a13][b369][m369];
        end
    endgenerate
    generate 
        localparam integer b370 = 6;
        for (m370 = 0; m370 < 16; m370 = m370 + 1) 
        begin: inbit370
            assign data_11[m370 + b370*16 + a13*28*16] = data_11_array[a13][b370][m370];
        end
    endgenerate
    generate 
        localparam integer b371 = 7;
        for (m371 = 0; m371 < 16; m371 = m371 + 1) 
        begin: inbit371
            assign data_11[m371 + b371*16 + a13*28*16] = data_11_array[a13][b371][m371];
        end
    endgenerate
    generate 
        localparam integer b372 = 8;
        for (m372 = 0; m372 < 16; m372 = m372 + 1) 
        begin: inbit372
            assign data_11[m372 + b372*16 + a13*28*16] = data_11_array[a13][b372][m372];
        end
    endgenerate
    generate 
        localparam integer b373 = 9;
        for (m373 = 0; m373 < 16; m373 = m373 + 1) 
        begin: inbit373
            assign data_11[m373 + b373*16 + a13*28*16] = data_11_array[a13][b373][m373];
        end
    endgenerate
    generate 
        localparam integer b374 = 10;
        for (m374 = 0; m374 < 16; m374 = m374 + 1) 
        begin: inbit374
            assign data_11[m374 + b374*16 + a13*28*16] = data_11_array[a13][b374][m374];
        end
    endgenerate
    generate 
        localparam integer b375 = 11;
        for (m375 = 0; m375 < 16; m375 = m375 + 1) 
        begin: inbit375
            assign data_11[m375 + b375*16 + a13*28*16] = data_11_array[a13][b375][m375];
        end
    endgenerate
    generate 
        localparam integer b376 = 12;
        for (m376 = 0; m376 < 16; m376 = m376 + 1) 
        begin: inbit376
            assign data_11[m376 + b376*16 + a13*28*16] = data_11_array[a13][b376][m376];
        end
    endgenerate
    generate 
        localparam integer b377 = 13;
        for (m377 = 0; m377 < 16; m377 = m377 + 1) 
        begin: inbit377
            assign data_11[m377 + b377*16 + a13*28*16] = data_11_array[a13][b377][m377];
        end
    endgenerate
    generate 
        localparam integer b378 = 14;
        for (m378 = 0; m378 < 16; m378 = m378 + 1) 
        begin: inbit378
            assign data_11[m378 + b378*16 + a13*28*16] = data_11_array[a13][b378][m378];
        end
    endgenerate
    generate 
        localparam integer b379 = 15;
        for (m379 = 0; m379 < 16; m379 = m379 + 1) 
        begin: inbit379
            assign data_11[m379 + b379*16 + a13*28*16] = data_11_array[a13][b379][m379];
        end
    endgenerate
    generate 
        localparam integer b380 = 16;
        for (m380 = 0; m380 < 16; m380 = m380 + 1) 
        begin: inbit380
            assign data_11[m380 + b380*16 + a13*28*16] = data_11_array[a13][b380][m380];
        end
    endgenerate
    generate 
        localparam integer b381 = 17;
        for (m381 = 0; m381 < 16; m381 = m381 + 1) 
        begin: inbit381
            assign data_11[m381 + b381*16 + a13*28*16] = data_11_array[a13][b381][m381];
        end
    endgenerate
    generate 
        localparam integer b382 = 18;
        for (m382 = 0; m382 < 16; m382 = m382 + 1) 
        begin: inbit382
            assign data_11[m382 + b382*16 + a13*28*16] = data_11_array[a13][b382][m382];
        end
    endgenerate
    generate 
        localparam integer b383 = 19;
        for (m383 = 0; m383 < 16; m383 = m383 + 1) 
        begin: inbit383
            assign data_11[m383 + b383*16 + a13*28*16] = data_11_array[a13][b383][m383];
        end
    endgenerate
    generate 
        localparam integer b384 = 20;
        for (m384 = 0; m384 < 16; m384 = m384 + 1) 
        begin: inbit384
            assign data_11[m384 + b384*16 + a13*28*16] = data_11_array[a13][b384][m384];
        end
    endgenerate
    generate 
        localparam integer b385 = 21;
        for (m385 = 0; m385 < 16; m385 = m385 + 1) 
        begin: inbit385
            assign data_11[m385 + b385*16 + a13*28*16] = data_11_array[a13][b385][m385];
        end
    endgenerate
    generate 
        localparam integer b386 = 22;
        for (m386 = 0; m386 < 16; m386 = m386 + 1) 
        begin: inbit386
            assign data_11[m386 + b386*16 + a13*28*16] = data_11_array[a13][b386][m386];
        end
    endgenerate
    generate 
        localparam integer b387 = 23;
        for (m387 = 0; m387 < 16; m387 = m387 + 1) 
        begin: inbit387
            assign data_11[m387 + b387*16 + a13*28*16] = data_11_array[a13][b387][m387];
        end
    endgenerate
    generate 
        localparam integer b388 = 24;
        for (m388 = 0; m388 < 16; m388 = m388 + 1) 
        begin: inbit388
            assign data_11[m388 + b388*16 + a13*28*16] = data_11_array[a13][b388][m388];
        end
    endgenerate
    generate 
        localparam integer b389 = 25;
        for (m389 = 0; m389 < 16; m389 = m389 + 1) 
        begin: inbit389
            assign data_11[m389 + b389*16 + a13*28*16] = data_11_array[a13][b389][m389];
        end
    endgenerate
    generate 
        localparam integer b390 = 26;
        for (m390 = 0; m390 < 16; m390 = m390 + 1) 
        begin: inbit390
            assign data_11[m390 + b390*16 + a13*28*16] = data_11_array[a13][b390][m390];
        end
    endgenerate
    generate 
        localparam integer b391 = 27;
        for (m391 = 0; m391 < 16; m391 = m391 + 1) 
        begin: inbit391
            assign data_11[m391 + b391*16 + a13*28*16] = data_11_array[a13][b391][m391];
        end
    endgenerate
    localparam integer a14 = 14;
    generate 
        localparam integer b392 = 0;
        for (m392 = 0; m392 < 16; m392 = m392 + 1) 
        begin: inbit392
            assign data_11[m392 + b392*16 + a14*28*16] = data_11_array[a14][b392][m392];
        end
    endgenerate
    generate 
        localparam integer b393 = 1;
        for (m393 = 0; m393 < 16; m393 = m393 + 1) 
        begin: inbit393
            assign data_11[m393 + b393*16 + a14*28*16] = data_11_array[a14][b393][m393];
        end
    endgenerate
    generate 
        localparam integer b394 = 2;
        for (m394 = 0; m394 < 16; m394 = m394 + 1) 
        begin: inbit394
            assign data_11[m394 + b394*16 + a14*28*16] = data_11_array[a14][b394][m394];
        end
    endgenerate
    generate 
        localparam integer b395 = 3;
        for (m395 = 0; m395 < 16; m395 = m395 + 1) 
        begin: inbit395
            assign data_11[m395 + b395*16 + a14*28*16] = data_11_array[a14][b395][m395];
        end
    endgenerate
    generate 
        localparam integer b396 = 4;
        for (m396 = 0; m396 < 16; m396 = m396 + 1) 
        begin: inbit396
            assign data_11[m396 + b396*16 + a14*28*16] = data_11_array[a14][b396][m396];
        end
    endgenerate
    generate 
        localparam integer b397 = 5;
        for (m397 = 0; m397 < 16; m397 = m397 + 1) 
        begin: inbit397
            assign data_11[m397 + b397*16 + a14*28*16] = data_11_array[a14][b397][m397];
        end
    endgenerate
    generate 
        localparam integer b398 = 6;
        for (m398 = 0; m398 < 16; m398 = m398 + 1) 
        begin: inbit398
            assign data_11[m398 + b398*16 + a14*28*16] = data_11_array[a14][b398][m398];
        end
    endgenerate
    generate 
        localparam integer b399 = 7;
        for (m399 = 0; m399 < 16; m399 = m399 + 1) 
        begin: inbit399
            assign data_11[m399 + b399*16 + a14*28*16] = data_11_array[a14][b399][m399];
        end
    endgenerate
    generate 
        localparam integer b400 = 8;
        for (m400 = 0; m400 < 16; m400 = m400 + 1) 
        begin: inbit400
            assign data_11[m400 + b400*16 + a14*28*16] = data_11_array[a14][b400][m400];
        end
    endgenerate
    generate 
        localparam integer b401 = 9;
        for (m401 = 0; m401 < 16; m401 = m401 + 1) 
        begin: inbit401
            assign data_11[m401 + b401*16 + a14*28*16] = data_11_array[a14][b401][m401];
        end
    endgenerate
    generate 
        localparam integer b402 = 10;
        for (m402 = 0; m402 < 16; m402 = m402 + 1) 
        begin: inbit402
            assign data_11[m402 + b402*16 + a14*28*16] = data_11_array[a14][b402][m402];
        end
    endgenerate
    generate 
        localparam integer b403 = 11;
        for (m403 = 0; m403 < 16; m403 = m403 + 1) 
        begin: inbit403
            assign data_11[m403 + b403*16 + a14*28*16] = data_11_array[a14][b403][m403];
        end
    endgenerate
    generate 
        localparam integer b404 = 12;
        for (m404 = 0; m404 < 16; m404 = m404 + 1) 
        begin: inbit404
            assign data_11[m404 + b404*16 + a14*28*16] = data_11_array[a14][b404][m404];
        end
    endgenerate
    generate 
        localparam integer b405 = 13;
        for (m405 = 0; m405 < 16; m405 = m405 + 1) 
        begin: inbit405
            assign data_11[m405 + b405*16 + a14*28*16] = data_11_array[a14][b405][m405];
        end
    endgenerate
    generate 
        localparam integer b406 = 14;
        for (m406 = 0; m406 < 16; m406 = m406 + 1) 
        begin: inbit406
            assign data_11[m406 + b406*16 + a14*28*16] = data_11_array[a14][b406][m406];
        end
    endgenerate
    generate 
        localparam integer b407 = 15;
        for (m407 = 0; m407 < 16; m407 = m407 + 1) 
        begin: inbit407
            assign data_11[m407 + b407*16 + a14*28*16] = data_11_array[a14][b407][m407];
        end
    endgenerate
    generate 
        localparam integer b408 = 16;
        for (m408 = 0; m408 < 16; m408 = m408 + 1) 
        begin: inbit408
            assign data_11[m408 + b408*16 + a14*28*16] = data_11_array[a14][b408][m408];
        end
    endgenerate
    generate 
        localparam integer b409 = 17;
        for (m409 = 0; m409 < 16; m409 = m409 + 1) 
        begin: inbit409
            assign data_11[m409 + b409*16 + a14*28*16] = data_11_array[a14][b409][m409];
        end
    endgenerate
    generate 
        localparam integer b410 = 18;
        for (m410 = 0; m410 < 16; m410 = m410 + 1) 
        begin: inbit410
            assign data_11[m410 + b410*16 + a14*28*16] = data_11_array[a14][b410][m410];
        end
    endgenerate
    generate 
        localparam integer b411 = 19;
        for (m411 = 0; m411 < 16; m411 = m411 + 1) 
        begin: inbit411
            assign data_11[m411 + b411*16 + a14*28*16] = data_11_array[a14][b411][m411];
        end
    endgenerate
    generate 
        localparam integer b412 = 20;
        for (m412 = 0; m412 < 16; m412 = m412 + 1) 
        begin: inbit412
            assign data_11[m412 + b412*16 + a14*28*16] = data_11_array[a14][b412][m412];
        end
    endgenerate
    generate 
        localparam integer b413 = 21;
        for (m413 = 0; m413 < 16; m413 = m413 + 1) 
        begin: inbit413
            assign data_11[m413 + b413*16 + a14*28*16] = data_11_array[a14][b413][m413];
        end
    endgenerate
    generate 
        localparam integer b414 = 22;
        for (m414 = 0; m414 < 16; m414 = m414 + 1) 
        begin: inbit414
            assign data_11[m414 + b414*16 + a14*28*16] = data_11_array[a14][b414][m414];
        end
    endgenerate
    generate 
        localparam integer b415 = 23;
        for (m415 = 0; m415 < 16; m415 = m415 + 1) 
        begin: inbit415
            assign data_11[m415 + b415*16 + a14*28*16] = data_11_array[a14][b415][m415];
        end
    endgenerate
    generate 
        localparam integer b416 = 24;
        for (m416 = 0; m416 < 16; m416 = m416 + 1) 
        begin: inbit416
            assign data_11[m416 + b416*16 + a14*28*16] = data_11_array[a14][b416][m416];
        end
    endgenerate
    generate 
        localparam integer b417 = 25;
        for (m417 = 0; m417 < 16; m417 = m417 + 1) 
        begin: inbit417
            assign data_11[m417 + b417*16 + a14*28*16] = data_11_array[a14][b417][m417];
        end
    endgenerate
    generate 
        localparam integer b418 = 26;
        for (m418 = 0; m418 < 16; m418 = m418 + 1) 
        begin: inbit418
            assign data_11[m418 + b418*16 + a14*28*16] = data_11_array[a14][b418][m418];
        end
    endgenerate
    generate 
        localparam integer b419 = 27;
        for (m419 = 0; m419 < 16; m419 = m419 + 1) 
        begin: inbit419
            assign data_11[m419 + b419*16 + a14*28*16] = data_11_array[a14][b419][m419];
        end
    endgenerate
    localparam integer a15 = 15;
    generate 
        localparam integer b420 = 0;
        for (m420 = 0; m420 < 16; m420 = m420 + 1) 
        begin: inbit420
            assign data_11[m420 + b420*16 + a15*28*16] = data_11_array[a15][b420][m420];
        end
    endgenerate
    generate 
        localparam integer b421 = 1;
        for (m421 = 0; m421 < 16; m421 = m421 + 1) 
        begin: inbit421
            assign data_11[m421 + b421*16 + a15*28*16] = data_11_array[a15][b421][m421];
        end
    endgenerate
    generate 
        localparam integer b422 = 2;
        for (m422 = 0; m422 < 16; m422 = m422 + 1) 
        begin: inbit422
            assign data_11[m422 + b422*16 + a15*28*16] = data_11_array[a15][b422][m422];
        end
    endgenerate
    generate 
        localparam integer b423 = 3;
        for (m423 = 0; m423 < 16; m423 = m423 + 1) 
        begin: inbit423
            assign data_11[m423 + b423*16 + a15*28*16] = data_11_array[a15][b423][m423];
        end
    endgenerate
    generate 
        localparam integer b424 = 4;
        for (m424 = 0; m424 < 16; m424 = m424 + 1) 
        begin: inbit424
            assign data_11[m424 + b424*16 + a15*28*16] = data_11_array[a15][b424][m424];
        end
    endgenerate
    generate 
        localparam integer b425 = 5;
        for (m425 = 0; m425 < 16; m425 = m425 + 1) 
        begin: inbit425
            assign data_11[m425 + b425*16 + a15*28*16] = data_11_array[a15][b425][m425];
        end
    endgenerate
    generate 
        localparam integer b426 = 6;
        for (m426 = 0; m426 < 16; m426 = m426 + 1) 
        begin: inbit426
            assign data_11[m426 + b426*16 + a15*28*16] = data_11_array[a15][b426][m426];
        end
    endgenerate
    generate 
        localparam integer b427 = 7;
        for (m427 = 0; m427 < 16; m427 = m427 + 1) 
        begin: inbit427
            assign data_11[m427 + b427*16 + a15*28*16] = data_11_array[a15][b427][m427];
        end
    endgenerate
    generate 
        localparam integer b428 = 8;
        for (m428 = 0; m428 < 16; m428 = m428 + 1) 
        begin: inbit428
            assign data_11[m428 + b428*16 + a15*28*16] = data_11_array[a15][b428][m428];
        end
    endgenerate
    generate 
        localparam integer b429 = 9;
        for (m429 = 0; m429 < 16; m429 = m429 + 1) 
        begin: inbit429
            assign data_11[m429 + b429*16 + a15*28*16] = data_11_array[a15][b429][m429];
        end
    endgenerate
    generate 
        localparam integer b430 = 10;
        for (m430 = 0; m430 < 16; m430 = m430 + 1) 
        begin: inbit430
            assign data_11[m430 + b430*16 + a15*28*16] = data_11_array[a15][b430][m430];
        end
    endgenerate
    generate 
        localparam integer b431 = 11;
        for (m431 = 0; m431 < 16; m431 = m431 + 1) 
        begin: inbit431
            assign data_11[m431 + b431*16 + a15*28*16] = data_11_array[a15][b431][m431];
        end
    endgenerate
    generate 
        localparam integer b432 = 12;
        for (m432 = 0; m432 < 16; m432 = m432 + 1) 
        begin: inbit432
            assign data_11[m432 + b432*16 + a15*28*16] = data_11_array[a15][b432][m432];
        end
    endgenerate
    generate 
        localparam integer b433 = 13;
        for (m433 = 0; m433 < 16; m433 = m433 + 1) 
        begin: inbit433
            assign data_11[m433 + b433*16 + a15*28*16] = data_11_array[a15][b433][m433];
        end
    endgenerate
    generate 
        localparam integer b434 = 14;
        for (m434 = 0; m434 < 16; m434 = m434 + 1) 
        begin: inbit434
            assign data_11[m434 + b434*16 + a15*28*16] = data_11_array[a15][b434][m434];
        end
    endgenerate
    generate 
        localparam integer b435 = 15;
        for (m435 = 0; m435 < 16; m435 = m435 + 1) 
        begin: inbit435
            assign data_11[m435 + b435*16 + a15*28*16] = data_11_array[a15][b435][m435];
        end
    endgenerate
    generate 
        localparam integer b436 = 16;
        for (m436 = 0; m436 < 16; m436 = m436 + 1) 
        begin: inbit436
            assign data_11[m436 + b436*16 + a15*28*16] = data_11_array[a15][b436][m436];
        end
    endgenerate
    generate 
        localparam integer b437 = 17;
        for (m437 = 0; m437 < 16; m437 = m437 + 1) 
        begin: inbit437
            assign data_11[m437 + b437*16 + a15*28*16] = data_11_array[a15][b437][m437];
        end
    endgenerate
    generate 
        localparam integer b438 = 18;
        for (m438 = 0; m438 < 16; m438 = m438 + 1) 
        begin: inbit438
            assign data_11[m438 + b438*16 + a15*28*16] = data_11_array[a15][b438][m438];
        end
    endgenerate
    generate 
        localparam integer b439 = 19;
        for (m439 = 0; m439 < 16; m439 = m439 + 1) 
        begin: inbit439
            assign data_11[m439 + b439*16 + a15*28*16] = data_11_array[a15][b439][m439];
        end
    endgenerate
    generate 
        localparam integer b440 = 20;
        for (m440 = 0; m440 < 16; m440 = m440 + 1) 
        begin: inbit440
            assign data_11[m440 + b440*16 + a15*28*16] = data_11_array[a15][b440][m440];
        end
    endgenerate
    generate 
        localparam integer b441 = 21;
        for (m441 = 0; m441 < 16; m441 = m441 + 1) 
        begin: inbit441
            assign data_11[m441 + b441*16 + a15*28*16] = data_11_array[a15][b441][m441];
        end
    endgenerate
    generate 
        localparam integer b442 = 22;
        for (m442 = 0; m442 < 16; m442 = m442 + 1) 
        begin: inbit442
            assign data_11[m442 + b442*16 + a15*28*16] = data_11_array[a15][b442][m442];
        end
    endgenerate
    generate 
        localparam integer b443 = 23;
        for (m443 = 0; m443 < 16; m443 = m443 + 1) 
        begin: inbit443
            assign data_11[m443 + b443*16 + a15*28*16] = data_11_array[a15][b443][m443];
        end
    endgenerate
    generate 
        localparam integer b444 = 24;
        for (m444 = 0; m444 < 16; m444 = m444 + 1) 
        begin: inbit444
            assign data_11[m444 + b444*16 + a15*28*16] = data_11_array[a15][b444][m444];
        end
    endgenerate
    generate 
        localparam integer b445 = 25;
        for (m445 = 0; m445 < 16; m445 = m445 + 1) 
        begin: inbit445
            assign data_11[m445 + b445*16 + a15*28*16] = data_11_array[a15][b445][m445];
        end
    endgenerate
    generate 
        localparam integer b446 = 26;
        for (m446 = 0; m446 < 16; m446 = m446 + 1) 
        begin: inbit446
            assign data_11[m446 + b446*16 + a15*28*16] = data_11_array[a15][b446][m446];
        end
    endgenerate
    generate 
        localparam integer b447 = 27;
        for (m447 = 0; m447 < 16; m447 = m447 + 1) 
        begin: inbit447
            assign data_11[m447 + b447*16 + a15*28*16] = data_11_array[a15][b447][m447];
        end
    endgenerate
    localparam integer a16 = 16;
    generate 
        localparam integer b448 = 0;
        for (m448 = 0; m448 < 16; m448 = m448 + 1) 
        begin: inbit448
            assign data_11[m448 + b448*16 + a16*28*16] = data_11_array[a16][b448][m448];
        end
    endgenerate
    generate 
        localparam integer b449 = 1;
        for (m449 = 0; m449 < 16; m449 = m449 + 1) 
        begin: inbit449
            assign data_11[m449 + b449*16 + a16*28*16] = data_11_array[a16][b449][m449];
        end
    endgenerate
    generate 
        localparam integer b450 = 2;
        for (m450 = 0; m450 < 16; m450 = m450 + 1) 
        begin: inbit450
            assign data_11[m450 + b450*16 + a16*28*16] = data_11_array[a16][b450][m450];
        end
    endgenerate
    generate 
        localparam integer b451 = 3;
        for (m451 = 0; m451 < 16; m451 = m451 + 1) 
        begin: inbit451
            assign data_11[m451 + b451*16 + a16*28*16] = data_11_array[a16][b451][m451];
        end
    endgenerate
    generate 
        localparam integer b452 = 4;
        for (m452 = 0; m452 < 16; m452 = m452 + 1) 
        begin: inbit452
            assign data_11[m452 + b452*16 + a16*28*16] = data_11_array[a16][b452][m452];
        end
    endgenerate
    generate 
        localparam integer b453 = 5;
        for (m453 = 0; m453 < 16; m453 = m453 + 1) 
        begin: inbit453
            assign data_11[m453 + b453*16 + a16*28*16] = data_11_array[a16][b453][m453];
        end
    endgenerate
    generate 
        localparam integer b454 = 6;
        for (m454 = 0; m454 < 16; m454 = m454 + 1) 
        begin: inbit454
            assign data_11[m454 + b454*16 + a16*28*16] = data_11_array[a16][b454][m454];
        end
    endgenerate
    generate 
        localparam integer b455 = 7;
        for (m455 = 0; m455 < 16; m455 = m455 + 1) 
        begin: inbit455
            assign data_11[m455 + b455*16 + a16*28*16] = data_11_array[a16][b455][m455];
        end
    endgenerate
    generate 
        localparam integer b456 = 8;
        for (m456 = 0; m456 < 16; m456 = m456 + 1) 
        begin: inbit456
            assign data_11[m456 + b456*16 + a16*28*16] = data_11_array[a16][b456][m456];
        end
    endgenerate
    generate 
        localparam integer b457 = 9;
        for (m457 = 0; m457 < 16; m457 = m457 + 1) 
        begin: inbit457
            assign data_11[m457 + b457*16 + a16*28*16] = data_11_array[a16][b457][m457];
        end
    endgenerate
    generate 
        localparam integer b458 = 10;
        for (m458 = 0; m458 < 16; m458 = m458 + 1) 
        begin: inbit458
            assign data_11[m458 + b458*16 + a16*28*16] = data_11_array[a16][b458][m458];
        end
    endgenerate
    generate 
        localparam integer b459 = 11;
        for (m459 = 0; m459 < 16; m459 = m459 + 1) 
        begin: inbit459
            assign data_11[m459 + b459*16 + a16*28*16] = data_11_array[a16][b459][m459];
        end
    endgenerate
    generate 
        localparam integer b460 = 12;
        for (m460 = 0; m460 < 16; m460 = m460 + 1) 
        begin: inbit460
            assign data_11[m460 + b460*16 + a16*28*16] = data_11_array[a16][b460][m460];
        end
    endgenerate
    generate 
        localparam integer b461 = 13;
        for (m461 = 0; m461 < 16; m461 = m461 + 1) 
        begin: inbit461
            assign data_11[m461 + b461*16 + a16*28*16] = data_11_array[a16][b461][m461];
        end
    endgenerate
    generate 
        localparam integer b462 = 14;
        for (m462 = 0; m462 < 16; m462 = m462 + 1) 
        begin: inbit462
            assign data_11[m462 + b462*16 + a16*28*16] = data_11_array[a16][b462][m462];
        end
    endgenerate
    generate 
        localparam integer b463 = 15;
        for (m463 = 0; m463 < 16; m463 = m463 + 1) 
        begin: inbit463
            assign data_11[m463 + b463*16 + a16*28*16] = data_11_array[a16][b463][m463];
        end
    endgenerate
    generate 
        localparam integer b464 = 16;
        for (m464 = 0; m464 < 16; m464 = m464 + 1) 
        begin: inbit464
            assign data_11[m464 + b464*16 + a16*28*16] = data_11_array[a16][b464][m464];
        end
    endgenerate
    generate 
        localparam integer b465 = 17;
        for (m465 = 0; m465 < 16; m465 = m465 + 1) 
        begin: inbit465
            assign data_11[m465 + b465*16 + a16*28*16] = data_11_array[a16][b465][m465];
        end
    endgenerate
    generate 
        localparam integer b466 = 18;
        for (m466 = 0; m466 < 16; m466 = m466 + 1) 
        begin: inbit466
            assign data_11[m466 + b466*16 + a16*28*16] = data_11_array[a16][b466][m466];
        end
    endgenerate
    generate 
        localparam integer b467 = 19;
        for (m467 = 0; m467 < 16; m467 = m467 + 1) 
        begin: inbit467
            assign data_11[m467 + b467*16 + a16*28*16] = data_11_array[a16][b467][m467];
        end
    endgenerate
    generate 
        localparam integer b468 = 20;
        for (m468 = 0; m468 < 16; m468 = m468 + 1) 
        begin: inbit468
            assign data_11[m468 + b468*16 + a16*28*16] = data_11_array[a16][b468][m468];
        end
    endgenerate
    generate 
        localparam integer b469 = 21;
        for (m469 = 0; m469 < 16; m469 = m469 + 1) 
        begin: inbit469
            assign data_11[m469 + b469*16 + a16*28*16] = data_11_array[a16][b469][m469];
        end
    endgenerate
    generate 
        localparam integer b470 = 22;
        for (m470 = 0; m470 < 16; m470 = m470 + 1) 
        begin: inbit470
            assign data_11[m470 + b470*16 + a16*28*16] = data_11_array[a16][b470][m470];
        end
    endgenerate
    generate 
        localparam integer b471 = 23;
        for (m471 = 0; m471 < 16; m471 = m471 + 1) 
        begin: inbit471
            assign data_11[m471 + b471*16 + a16*28*16] = data_11_array[a16][b471][m471];
        end
    endgenerate
    generate 
        localparam integer b472 = 24;
        for (m472 = 0; m472 < 16; m472 = m472 + 1) 
        begin: inbit472
            assign data_11[m472 + b472*16 + a16*28*16] = data_11_array[a16][b472][m472];
        end
    endgenerate
    generate 
        localparam integer b473 = 25;
        for (m473 = 0; m473 < 16; m473 = m473 + 1) 
        begin: inbit473
            assign data_11[m473 + b473*16 + a16*28*16] = data_11_array[a16][b473][m473];
        end
    endgenerate
    generate 
        localparam integer b474 = 26;
        for (m474 = 0; m474 < 16; m474 = m474 + 1) 
        begin: inbit474
            assign data_11[m474 + b474*16 + a16*28*16] = data_11_array[a16][b474][m474];
        end
    endgenerate
    generate 
        localparam integer b475 = 27;
        for (m475 = 0; m475 < 16; m475 = m475 + 1) 
        begin: inbit475
            assign data_11[m475 + b475*16 + a16*28*16] = data_11_array[a16][b475][m475];
        end
    endgenerate
    localparam integer a17 = 17;
    generate 
        localparam integer b476 = 0;
        for (m476 = 0; m476 < 16; m476 = m476 + 1) 
        begin: inbit476
            assign data_11[m476 + b476*16 + a17*28*16] = data_11_array[a17][b476][m476];
        end
    endgenerate
    generate 
        localparam integer b477 = 1;
        for (m477 = 0; m477 < 16; m477 = m477 + 1) 
        begin: inbit477
            assign data_11[m477 + b477*16 + a17*28*16] = data_11_array[a17][b477][m477];
        end
    endgenerate
    generate 
        localparam integer b478 = 2;
        for (m478 = 0; m478 < 16; m478 = m478 + 1) 
        begin: inbit478
            assign data_11[m478 + b478*16 + a17*28*16] = data_11_array[a17][b478][m478];
        end
    endgenerate
    generate 
        localparam integer b479 = 3;
        for (m479 = 0; m479 < 16; m479 = m479 + 1) 
        begin: inbit479
            assign data_11[m479 + b479*16 + a17*28*16] = data_11_array[a17][b479][m479];
        end
    endgenerate
    generate 
        localparam integer b480 = 4;
        for (m480 = 0; m480 < 16; m480 = m480 + 1) 
        begin: inbit480
            assign data_11[m480 + b480*16 + a17*28*16] = data_11_array[a17][b480][m480];
        end
    endgenerate
    generate 
        localparam integer b481 = 5;
        for (m481 = 0; m481 < 16; m481 = m481 + 1) 
        begin: inbit481
            assign data_11[m481 + b481*16 + a17*28*16] = data_11_array[a17][b481][m481];
        end
    endgenerate
    generate 
        localparam integer b482 = 6;
        for (m482 = 0; m482 < 16; m482 = m482 + 1) 
        begin: inbit482
            assign data_11[m482 + b482*16 + a17*28*16] = data_11_array[a17][b482][m482];
        end
    endgenerate
    generate 
        localparam integer b483 = 7;
        for (m483 = 0; m483 < 16; m483 = m483 + 1) 
        begin: inbit483
            assign data_11[m483 + b483*16 + a17*28*16] = data_11_array[a17][b483][m483];
        end
    endgenerate
    generate 
        localparam integer b484 = 8;
        for (m484 = 0; m484 < 16; m484 = m484 + 1) 
        begin: inbit484
            assign data_11[m484 + b484*16 + a17*28*16] = data_11_array[a17][b484][m484];
        end
    endgenerate
    generate 
        localparam integer b485 = 9;
        for (m485 = 0; m485 < 16; m485 = m485 + 1) 
        begin: inbit485
            assign data_11[m485 + b485*16 + a17*28*16] = data_11_array[a17][b485][m485];
        end
    endgenerate
    generate 
        localparam integer b486 = 10;
        for (m486 = 0; m486 < 16; m486 = m486 + 1) 
        begin: inbit486
            assign data_11[m486 + b486*16 + a17*28*16] = data_11_array[a17][b486][m486];
        end
    endgenerate
    generate 
        localparam integer b487 = 11;
        for (m487 = 0; m487 < 16; m487 = m487 + 1) 
        begin: inbit487
            assign data_11[m487 + b487*16 + a17*28*16] = data_11_array[a17][b487][m487];
        end
    endgenerate
    generate 
        localparam integer b488 = 12;
        for (m488 = 0; m488 < 16; m488 = m488 + 1) 
        begin: inbit488
            assign data_11[m488 + b488*16 + a17*28*16] = data_11_array[a17][b488][m488];
        end
    endgenerate
    generate 
        localparam integer b489 = 13;
        for (m489 = 0; m489 < 16; m489 = m489 + 1) 
        begin: inbit489
            assign data_11[m489 + b489*16 + a17*28*16] = data_11_array[a17][b489][m489];
        end
    endgenerate
    generate 
        localparam integer b490 = 14;
        for (m490 = 0; m490 < 16; m490 = m490 + 1) 
        begin: inbit490
            assign data_11[m490 + b490*16 + a17*28*16] = data_11_array[a17][b490][m490];
        end
    endgenerate
    generate 
        localparam integer b491 = 15;
        for (m491 = 0; m491 < 16; m491 = m491 + 1) 
        begin: inbit491
            assign data_11[m491 + b491*16 + a17*28*16] = data_11_array[a17][b491][m491];
        end
    endgenerate
    generate 
        localparam integer b492 = 16;
        for (m492 = 0; m492 < 16; m492 = m492 + 1) 
        begin: inbit492
            assign data_11[m492 + b492*16 + a17*28*16] = data_11_array[a17][b492][m492];
        end
    endgenerate
    generate 
        localparam integer b493 = 17;
        for (m493 = 0; m493 < 16; m493 = m493 + 1) 
        begin: inbit493
            assign data_11[m493 + b493*16 + a17*28*16] = data_11_array[a17][b493][m493];
        end
    endgenerate
    generate 
        localparam integer b494 = 18;
        for (m494 = 0; m494 < 16; m494 = m494 + 1) 
        begin: inbit494
            assign data_11[m494 + b494*16 + a17*28*16] = data_11_array[a17][b494][m494];
        end
    endgenerate
    generate 
        localparam integer b495 = 19;
        for (m495 = 0; m495 < 16; m495 = m495 + 1) 
        begin: inbit495
            assign data_11[m495 + b495*16 + a17*28*16] = data_11_array[a17][b495][m495];
        end
    endgenerate
    generate 
        localparam integer b496 = 20;
        for (m496 = 0; m496 < 16; m496 = m496 + 1) 
        begin: inbit496
            assign data_11[m496 + b496*16 + a17*28*16] = data_11_array[a17][b496][m496];
        end
    endgenerate
    generate 
        localparam integer b497 = 21;
        for (m497 = 0; m497 < 16; m497 = m497 + 1) 
        begin: inbit497
            assign data_11[m497 + b497*16 + a17*28*16] = data_11_array[a17][b497][m497];
        end
    endgenerate
    generate 
        localparam integer b498 = 22;
        for (m498 = 0; m498 < 16; m498 = m498 + 1) 
        begin: inbit498
            assign data_11[m498 + b498*16 + a17*28*16] = data_11_array[a17][b498][m498];
        end
    endgenerate
    generate 
        localparam integer b499 = 23;
        for (m499 = 0; m499 < 16; m499 = m499 + 1) 
        begin: inbit499
            assign data_11[m499 + b499*16 + a17*28*16] = data_11_array[a17][b499][m499];
        end
    endgenerate
    generate 
        localparam integer b500 = 24;
        for (m500 = 0; m500 < 16; m500 = m500 + 1) 
        begin: inbit500
            assign data_11[m500 + b500*16 + a17*28*16] = data_11_array[a17][b500][m500];
        end
    endgenerate
    generate 
        localparam integer b501 = 25;
        for (m501 = 0; m501 < 16; m501 = m501 + 1) 
        begin: inbit501
            assign data_11[m501 + b501*16 + a17*28*16] = data_11_array[a17][b501][m501];
        end
    endgenerate
    generate 
        localparam integer b502 = 26;
        for (m502 = 0; m502 < 16; m502 = m502 + 1) 
        begin: inbit502
            assign data_11[m502 + b502*16 + a17*28*16] = data_11_array[a17][b502][m502];
        end
    endgenerate
    generate 
        localparam integer b503 = 27;
        for (m503 = 0; m503 < 16; m503 = m503 + 1) 
        begin: inbit503
            assign data_11[m503 + b503*16 + a17*28*16] = data_11_array[a17][b503][m503];
        end
    endgenerate
    localparam integer a18 = 18;
    generate 
        localparam integer b504 = 0;
        for (m504 = 0; m504 < 16; m504 = m504 + 1) 
        begin: inbit504
            assign data_11[m504 + b504*16 + a18*28*16] = data_11_array[a18][b504][m504];
        end
    endgenerate
    generate 
        localparam integer b505 = 1;
        for (m505 = 0; m505 < 16; m505 = m505 + 1) 
        begin: inbit505
            assign data_11[m505 + b505*16 + a18*28*16] = data_11_array[a18][b505][m505];
        end
    endgenerate
    generate 
        localparam integer b506 = 2;
        for (m506 = 0; m506 < 16; m506 = m506 + 1) 
        begin: inbit506
            assign data_11[m506 + b506*16 + a18*28*16] = data_11_array[a18][b506][m506];
        end
    endgenerate
    generate 
        localparam integer b507 = 3;
        for (m507 = 0; m507 < 16; m507 = m507 + 1) 
        begin: inbit507
            assign data_11[m507 + b507*16 + a18*28*16] = data_11_array[a18][b507][m507];
        end
    endgenerate
    generate 
        localparam integer b508 = 4;
        for (m508 = 0; m508 < 16; m508 = m508 + 1) 
        begin: inbit508
            assign data_11[m508 + b508*16 + a18*28*16] = data_11_array[a18][b508][m508];
        end
    endgenerate
    generate 
        localparam integer b509 = 5;
        for (m509 = 0; m509 < 16; m509 = m509 + 1) 
        begin: inbit509
            assign data_11[m509 + b509*16 + a18*28*16] = data_11_array[a18][b509][m509];
        end
    endgenerate
    generate 
        localparam integer b510 = 6;
        for (m510 = 0; m510 < 16; m510 = m510 + 1) 
        begin: inbit510
            assign data_11[m510 + b510*16 + a18*28*16] = data_11_array[a18][b510][m510];
        end
    endgenerate
    generate 
        localparam integer b511 = 7;
        for (m511 = 0; m511 < 16; m511 = m511 + 1) 
        begin: inbit511
            assign data_11[m511 + b511*16 + a18*28*16] = data_11_array[a18][b511][m511];
        end
    endgenerate
    generate 
        localparam integer b512 = 8;
        for (m512 = 0; m512 < 16; m512 = m512 + 1) 
        begin: inbit512
            assign data_11[m512 + b512*16 + a18*28*16] = data_11_array[a18][b512][m512];
        end
    endgenerate
    generate 
        localparam integer b513 = 9;
        for (m513 = 0; m513 < 16; m513 = m513 + 1) 
        begin: inbit513
            assign data_11[m513 + b513*16 + a18*28*16] = data_11_array[a18][b513][m513];
        end
    endgenerate
    generate 
        localparam integer b514 = 10;
        for (m514 = 0; m514 < 16; m514 = m514 + 1) 
        begin: inbit514
            assign data_11[m514 + b514*16 + a18*28*16] = data_11_array[a18][b514][m514];
        end
    endgenerate
    generate 
        localparam integer b515 = 11;
        for (m515 = 0; m515 < 16; m515 = m515 + 1) 
        begin: inbit515
            assign data_11[m515 + b515*16 + a18*28*16] = data_11_array[a18][b515][m515];
        end
    endgenerate
    generate 
        localparam integer b516 = 12;
        for (m516 = 0; m516 < 16; m516 = m516 + 1) 
        begin: inbit516
            assign data_11[m516 + b516*16 + a18*28*16] = data_11_array[a18][b516][m516];
        end
    endgenerate
    generate 
        localparam integer b517 = 13;
        for (m517 = 0; m517 < 16; m517 = m517 + 1) 
        begin: inbit517
            assign data_11[m517 + b517*16 + a18*28*16] = data_11_array[a18][b517][m517];
        end
    endgenerate
    generate 
        localparam integer b518 = 14;
        for (m518 = 0; m518 < 16; m518 = m518 + 1) 
        begin: inbit518
            assign data_11[m518 + b518*16 + a18*28*16] = data_11_array[a18][b518][m518];
        end
    endgenerate
    generate 
        localparam integer b519 = 15;
        for (m519 = 0; m519 < 16; m519 = m519 + 1) 
        begin: inbit519
            assign data_11[m519 + b519*16 + a18*28*16] = data_11_array[a18][b519][m519];
        end
    endgenerate
    generate 
        localparam integer b520 = 16;
        for (m520 = 0; m520 < 16; m520 = m520 + 1) 
        begin: inbit520
            assign data_11[m520 + b520*16 + a18*28*16] = data_11_array[a18][b520][m520];
        end
    endgenerate
    generate 
        localparam integer b521 = 17;
        for (m521 = 0; m521 < 16; m521 = m521 + 1) 
        begin: inbit521
            assign data_11[m521 + b521*16 + a18*28*16] = data_11_array[a18][b521][m521];
        end
    endgenerate
    generate 
        localparam integer b522 = 18;
        for (m522 = 0; m522 < 16; m522 = m522 + 1) 
        begin: inbit522
            assign data_11[m522 + b522*16 + a18*28*16] = data_11_array[a18][b522][m522];
        end
    endgenerate
    generate 
        localparam integer b523 = 19;
        for (m523 = 0; m523 < 16; m523 = m523 + 1) 
        begin: inbit523
            assign data_11[m523 + b523*16 + a18*28*16] = data_11_array[a18][b523][m523];
        end
    endgenerate
    generate 
        localparam integer b524 = 20;
        for (m524 = 0; m524 < 16; m524 = m524 + 1) 
        begin: inbit524
            assign data_11[m524 + b524*16 + a18*28*16] = data_11_array[a18][b524][m524];
        end
    endgenerate
    generate 
        localparam integer b525 = 21;
        for (m525 = 0; m525 < 16; m525 = m525 + 1) 
        begin: inbit525
            assign data_11[m525 + b525*16 + a18*28*16] = data_11_array[a18][b525][m525];
        end
    endgenerate
    generate 
        localparam integer b526 = 22;
        for (m526 = 0; m526 < 16; m526 = m526 + 1) 
        begin: inbit526
            assign data_11[m526 + b526*16 + a18*28*16] = data_11_array[a18][b526][m526];
        end
    endgenerate
    generate 
        localparam integer b527 = 23;
        for (m527 = 0; m527 < 16; m527 = m527 + 1) 
        begin: inbit527
            assign data_11[m527 + b527*16 + a18*28*16] = data_11_array[a18][b527][m527];
        end
    endgenerate
    generate 
        localparam integer b528 = 24;
        for (m528 = 0; m528 < 16; m528 = m528 + 1) 
        begin: inbit528
            assign data_11[m528 + b528*16 + a18*28*16] = data_11_array[a18][b528][m528];
        end
    endgenerate
    generate 
        localparam integer b529 = 25;
        for (m529 = 0; m529 < 16; m529 = m529 + 1) 
        begin: inbit529
            assign data_11[m529 + b529*16 + a18*28*16] = data_11_array[a18][b529][m529];
        end
    endgenerate
    generate 
        localparam integer b530 = 26;
        for (m530 = 0; m530 < 16; m530 = m530 + 1) 
        begin: inbit530
            assign data_11[m530 + b530*16 + a18*28*16] = data_11_array[a18][b530][m530];
        end
    endgenerate
    generate 
        localparam integer b531 = 27;
        for (m531 = 0; m531 < 16; m531 = m531 + 1) 
        begin: inbit531
            assign data_11[m531 + b531*16 + a18*28*16] = data_11_array[a18][b531][m531];
        end
    endgenerate
    localparam integer a19 = 19;
    generate 
        localparam integer b532 = 0;
        for (m532 = 0; m532 < 16; m532 = m532 + 1) 
        begin: inbit532
            assign data_11[m532 + b532*16 + a19*28*16] = data_11_array[a19][b532][m532];
        end
    endgenerate
    generate 
        localparam integer b533 = 1;
        for (m533 = 0; m533 < 16; m533 = m533 + 1) 
        begin: inbit533
            assign data_11[m533 + b533*16 + a19*28*16] = data_11_array[a19][b533][m533];
        end
    endgenerate
    generate 
        localparam integer b534 = 2;
        for (m534 = 0; m534 < 16; m534 = m534 + 1) 
        begin: inbit534
            assign data_11[m534 + b534*16 + a19*28*16] = data_11_array[a19][b534][m534];
        end
    endgenerate
    generate 
        localparam integer b535 = 3;
        for (m535 = 0; m535 < 16; m535 = m535 + 1) 
        begin: inbit535
            assign data_11[m535 + b535*16 + a19*28*16] = data_11_array[a19][b535][m535];
        end
    endgenerate
    generate 
        localparam integer b536 = 4;
        for (m536 = 0; m536 < 16; m536 = m536 + 1) 
        begin: inbit536
            assign data_11[m536 + b536*16 + a19*28*16] = data_11_array[a19][b536][m536];
        end
    endgenerate
    generate 
        localparam integer b537 = 5;
        for (m537 = 0; m537 < 16; m537 = m537 + 1) 
        begin: inbit537
            assign data_11[m537 + b537*16 + a19*28*16] = data_11_array[a19][b537][m537];
        end
    endgenerate
    generate 
        localparam integer b538 = 6;
        for (m538 = 0; m538 < 16; m538 = m538 + 1) 
        begin: inbit538
            assign data_11[m538 + b538*16 + a19*28*16] = data_11_array[a19][b538][m538];
        end
    endgenerate
    generate 
        localparam integer b539 = 7;
        for (m539 = 0; m539 < 16; m539 = m539 + 1) 
        begin: inbit539
            assign data_11[m539 + b539*16 + a19*28*16] = data_11_array[a19][b539][m539];
        end
    endgenerate
    generate 
        localparam integer b540 = 8;
        for (m540 = 0; m540 < 16; m540 = m540 + 1) 
        begin: inbit540
            assign data_11[m540 + b540*16 + a19*28*16] = data_11_array[a19][b540][m540];
        end
    endgenerate
    generate 
        localparam integer b541 = 9;
        for (m541 = 0; m541 < 16; m541 = m541 + 1) 
        begin: inbit541
            assign data_11[m541 + b541*16 + a19*28*16] = data_11_array[a19][b541][m541];
        end
    endgenerate
    generate 
        localparam integer b542 = 10;
        for (m542 = 0; m542 < 16; m542 = m542 + 1) 
        begin: inbit542
            assign data_11[m542 + b542*16 + a19*28*16] = data_11_array[a19][b542][m542];
        end
    endgenerate
    generate 
        localparam integer b543 = 11;
        for (m543 = 0; m543 < 16; m543 = m543 + 1) 
        begin: inbit543
            assign data_11[m543 + b543*16 + a19*28*16] = data_11_array[a19][b543][m543];
        end
    endgenerate
    generate 
        localparam integer b544 = 12;
        for (m544 = 0; m544 < 16; m544 = m544 + 1) 
        begin: inbit544
            assign data_11[m544 + b544*16 + a19*28*16] = data_11_array[a19][b544][m544];
        end
    endgenerate
    generate 
        localparam integer b545 = 13;
        for (m545 = 0; m545 < 16; m545 = m545 + 1) 
        begin: inbit545
            assign data_11[m545 + b545*16 + a19*28*16] = data_11_array[a19][b545][m545];
        end
    endgenerate
    generate 
        localparam integer b546 = 14;
        for (m546 = 0; m546 < 16; m546 = m546 + 1) 
        begin: inbit546
            assign data_11[m546 + b546*16 + a19*28*16] = data_11_array[a19][b546][m546];
        end
    endgenerate
    generate 
        localparam integer b547 = 15;
        for (m547 = 0; m547 < 16; m547 = m547 + 1) 
        begin: inbit547
            assign data_11[m547 + b547*16 + a19*28*16] = data_11_array[a19][b547][m547];
        end
    endgenerate
    generate 
        localparam integer b548 = 16;
        for (m548 = 0; m548 < 16; m548 = m548 + 1) 
        begin: inbit548
            assign data_11[m548 + b548*16 + a19*28*16] = data_11_array[a19][b548][m548];
        end
    endgenerate
    generate 
        localparam integer b549 = 17;
        for (m549 = 0; m549 < 16; m549 = m549 + 1) 
        begin: inbit549
            assign data_11[m549 + b549*16 + a19*28*16] = data_11_array[a19][b549][m549];
        end
    endgenerate
    generate 
        localparam integer b550 = 18;
        for (m550 = 0; m550 < 16; m550 = m550 + 1) 
        begin: inbit550
            assign data_11[m550 + b550*16 + a19*28*16] = data_11_array[a19][b550][m550];
        end
    endgenerate
    generate 
        localparam integer b551 = 19;
        for (m551 = 0; m551 < 16; m551 = m551 + 1) 
        begin: inbit551
            assign data_11[m551 + b551*16 + a19*28*16] = data_11_array[a19][b551][m551];
        end
    endgenerate
    generate 
        localparam integer b552 = 20;
        for (m552 = 0; m552 < 16; m552 = m552 + 1) 
        begin: inbit552
            assign data_11[m552 + b552*16 + a19*28*16] = data_11_array[a19][b552][m552];
        end
    endgenerate
    generate 
        localparam integer b553 = 21;
        for (m553 = 0; m553 < 16; m553 = m553 + 1) 
        begin: inbit553
            assign data_11[m553 + b553*16 + a19*28*16] = data_11_array[a19][b553][m553];
        end
    endgenerate
    generate 
        localparam integer b554 = 22;
        for (m554 = 0; m554 < 16; m554 = m554 + 1) 
        begin: inbit554
            assign data_11[m554 + b554*16 + a19*28*16] = data_11_array[a19][b554][m554];
        end
    endgenerate
    generate 
        localparam integer b555 = 23;
        for (m555 = 0; m555 < 16; m555 = m555 + 1) 
        begin: inbit555
            assign data_11[m555 + b555*16 + a19*28*16] = data_11_array[a19][b555][m555];
        end
    endgenerate
    generate 
        localparam integer b556 = 24;
        for (m556 = 0; m556 < 16; m556 = m556 + 1) 
        begin: inbit556
            assign data_11[m556 + b556*16 + a19*28*16] = data_11_array[a19][b556][m556];
        end
    endgenerate
    generate 
        localparam integer b557 = 25;
        for (m557 = 0; m557 < 16; m557 = m557 + 1) 
        begin: inbit557
            assign data_11[m557 + b557*16 + a19*28*16] = data_11_array[a19][b557][m557];
        end
    endgenerate
    generate 
        localparam integer b558 = 26;
        for (m558 = 0; m558 < 16; m558 = m558 + 1) 
        begin: inbit558
            assign data_11[m558 + b558*16 + a19*28*16] = data_11_array[a19][b558][m558];
        end
    endgenerate
    generate 
        localparam integer b559 = 27;
        for (m559 = 0; m559 < 16; m559 = m559 + 1) 
        begin: inbit559
            assign data_11[m559 + b559*16 + a19*28*16] = data_11_array[a19][b559][m559];
        end
    endgenerate
    localparam integer a20 = 20;
    generate 
        localparam integer b560 = 0;
        for (m560 = 0; m560 < 16; m560 = m560 + 1) 
        begin: inbit560
            assign data_11[m560 + b560*16 + a20*28*16] = data_11_array[a20][b560][m560];
        end
    endgenerate
    generate 
        localparam integer b561 = 1;
        for (m561 = 0; m561 < 16; m561 = m561 + 1) 
        begin: inbit561
            assign data_11[m561 + b561*16 + a20*28*16] = data_11_array[a20][b561][m561];
        end
    endgenerate
    generate 
        localparam integer b562 = 2;
        for (m562 = 0; m562 < 16; m562 = m562 + 1) 
        begin: inbit562
            assign data_11[m562 + b562*16 + a20*28*16] = data_11_array[a20][b562][m562];
        end
    endgenerate
    generate 
        localparam integer b563 = 3;
        for (m563 = 0; m563 < 16; m563 = m563 + 1) 
        begin: inbit563
            assign data_11[m563 + b563*16 + a20*28*16] = data_11_array[a20][b563][m563];
        end
    endgenerate
    generate 
        localparam integer b564 = 4;
        for (m564 = 0; m564 < 16; m564 = m564 + 1) 
        begin: inbit564
            assign data_11[m564 + b564*16 + a20*28*16] = data_11_array[a20][b564][m564];
        end
    endgenerate
    generate 
        localparam integer b565 = 5;
        for (m565 = 0; m565 < 16; m565 = m565 + 1) 
        begin: inbit565
            assign data_11[m565 + b565*16 + a20*28*16] = data_11_array[a20][b565][m565];
        end
    endgenerate
    generate 
        localparam integer b566 = 6;
        for (m566 = 0; m566 < 16; m566 = m566 + 1) 
        begin: inbit566
            assign data_11[m566 + b566*16 + a20*28*16] = data_11_array[a20][b566][m566];
        end
    endgenerate
    generate 
        localparam integer b567 = 7;
        for (m567 = 0; m567 < 16; m567 = m567 + 1) 
        begin: inbit567
            assign data_11[m567 + b567*16 + a20*28*16] = data_11_array[a20][b567][m567];
        end
    endgenerate
    generate 
        localparam integer b568 = 8;
        for (m568 = 0; m568 < 16; m568 = m568 + 1) 
        begin: inbit568
            assign data_11[m568 + b568*16 + a20*28*16] = data_11_array[a20][b568][m568];
        end
    endgenerate
    generate 
        localparam integer b569 = 9;
        for (m569 = 0; m569 < 16; m569 = m569 + 1) 
        begin: inbit569
            assign data_11[m569 + b569*16 + a20*28*16] = data_11_array[a20][b569][m569];
        end
    endgenerate
    generate 
        localparam integer b570 = 10;
        for (m570 = 0; m570 < 16; m570 = m570 + 1) 
        begin: inbit570
            assign data_11[m570 + b570*16 + a20*28*16] = data_11_array[a20][b570][m570];
        end
    endgenerate
    generate 
        localparam integer b571 = 11;
        for (m571 = 0; m571 < 16; m571 = m571 + 1) 
        begin: inbit571
            assign data_11[m571 + b571*16 + a20*28*16] = data_11_array[a20][b571][m571];
        end
    endgenerate
    generate 
        localparam integer b572 = 12;
        for (m572 = 0; m572 < 16; m572 = m572 + 1) 
        begin: inbit572
            assign data_11[m572 + b572*16 + a20*28*16] = data_11_array[a20][b572][m572];
        end
    endgenerate
    generate 
        localparam integer b573 = 13;
        for (m573 = 0; m573 < 16; m573 = m573 + 1) 
        begin: inbit573
            assign data_11[m573 + b573*16 + a20*28*16] = data_11_array[a20][b573][m573];
        end
    endgenerate
    generate 
        localparam integer b574 = 14;
        for (m574 = 0; m574 < 16; m574 = m574 + 1) 
        begin: inbit574
            assign data_11[m574 + b574*16 + a20*28*16] = data_11_array[a20][b574][m574];
        end
    endgenerate
    generate 
        localparam integer b575 = 15;
        for (m575 = 0; m575 < 16; m575 = m575 + 1) 
        begin: inbit575
            assign data_11[m575 + b575*16 + a20*28*16] = data_11_array[a20][b575][m575];
        end
    endgenerate
    generate 
        localparam integer b576 = 16;
        for (m576 = 0; m576 < 16; m576 = m576 + 1) 
        begin: inbit576
            assign data_11[m576 + b576*16 + a20*28*16] = data_11_array[a20][b576][m576];
        end
    endgenerate
    generate 
        localparam integer b577 = 17;
        for (m577 = 0; m577 < 16; m577 = m577 + 1) 
        begin: inbit577
            assign data_11[m577 + b577*16 + a20*28*16] = data_11_array[a20][b577][m577];
        end
    endgenerate
    generate 
        localparam integer b578 = 18;
        for (m578 = 0; m578 < 16; m578 = m578 + 1) 
        begin: inbit578
            assign data_11[m578 + b578*16 + a20*28*16] = data_11_array[a20][b578][m578];
        end
    endgenerate
    generate 
        localparam integer b579 = 19;
        for (m579 = 0; m579 < 16; m579 = m579 + 1) 
        begin: inbit579
            assign data_11[m579 + b579*16 + a20*28*16] = data_11_array[a20][b579][m579];
        end
    endgenerate
    generate 
        localparam integer b580 = 20;
        for (m580 = 0; m580 < 16; m580 = m580 + 1) 
        begin: inbit580
            assign data_11[m580 + b580*16 + a20*28*16] = data_11_array[a20][b580][m580];
        end
    endgenerate
    generate 
        localparam integer b581 = 21;
        for (m581 = 0; m581 < 16; m581 = m581 + 1) 
        begin: inbit581
            assign data_11[m581 + b581*16 + a20*28*16] = data_11_array[a20][b581][m581];
        end
    endgenerate
    generate 
        localparam integer b582 = 22;
        for (m582 = 0; m582 < 16; m582 = m582 + 1) 
        begin: inbit582
            assign data_11[m582 + b582*16 + a20*28*16] = data_11_array[a20][b582][m582];
        end
    endgenerate
    generate 
        localparam integer b583 = 23;
        for (m583 = 0; m583 < 16; m583 = m583 + 1) 
        begin: inbit583
            assign data_11[m583 + b583*16 + a20*28*16] = data_11_array[a20][b583][m583];
        end
    endgenerate
    generate 
        localparam integer b584 = 24;
        for (m584 = 0; m584 < 16; m584 = m584 + 1) 
        begin: inbit584
            assign data_11[m584 + b584*16 + a20*28*16] = data_11_array[a20][b584][m584];
        end
    endgenerate
    generate 
        localparam integer b585 = 25;
        for (m585 = 0; m585 < 16; m585 = m585 + 1) 
        begin: inbit585
            assign data_11[m585 + b585*16 + a20*28*16] = data_11_array[a20][b585][m585];
        end
    endgenerate
    generate 
        localparam integer b586 = 26;
        for (m586 = 0; m586 < 16; m586 = m586 + 1) 
        begin: inbit586
            assign data_11[m586 + b586*16 + a20*28*16] = data_11_array[a20][b586][m586];
        end
    endgenerate
    generate 
        localparam integer b587 = 27;
        for (m587 = 0; m587 < 16; m587 = m587 + 1) 
        begin: inbit587
            assign data_11[m587 + b587*16 + a20*28*16] = data_11_array[a20][b587][m587];
        end
    endgenerate
    localparam integer a21 = 21;
    generate 
        localparam integer b588 = 0;
        for (m588 = 0; m588 < 16; m588 = m588 + 1) 
        begin: inbit588
            assign data_11[m588 + b588*16 + a21*28*16] = data_11_array[a21][b588][m588];
        end
    endgenerate
    generate 
        localparam integer b589 = 1;
        for (m589 = 0; m589 < 16; m589 = m589 + 1) 
        begin: inbit589
            assign data_11[m589 + b589*16 + a21*28*16] = data_11_array[a21][b589][m589];
        end
    endgenerate
    generate 
        localparam integer b590 = 2;
        for (m590 = 0; m590 < 16; m590 = m590 + 1) 
        begin: inbit590
            assign data_11[m590 + b590*16 + a21*28*16] = data_11_array[a21][b590][m590];
        end
    endgenerate
    generate 
        localparam integer b591 = 3;
        for (m591 = 0; m591 < 16; m591 = m591 + 1) 
        begin: inbit591
            assign data_11[m591 + b591*16 + a21*28*16] = data_11_array[a21][b591][m591];
        end
    endgenerate
    generate 
        localparam integer b592 = 4;
        for (m592 = 0; m592 < 16; m592 = m592 + 1) 
        begin: inbit592
            assign data_11[m592 + b592*16 + a21*28*16] = data_11_array[a21][b592][m592];
        end
    endgenerate
    generate 
        localparam integer b593 = 5;
        for (m593 = 0; m593 < 16; m593 = m593 + 1) 
        begin: inbit593
            assign data_11[m593 + b593*16 + a21*28*16] = data_11_array[a21][b593][m593];
        end
    endgenerate
    generate 
        localparam integer b594 = 6;
        for (m594 = 0; m594 < 16; m594 = m594 + 1) 
        begin: inbit594
            assign data_11[m594 + b594*16 + a21*28*16] = data_11_array[a21][b594][m594];
        end
    endgenerate
    generate 
        localparam integer b595 = 7;
        for (m595 = 0; m595 < 16; m595 = m595 + 1) 
        begin: inbit595
            assign data_11[m595 + b595*16 + a21*28*16] = data_11_array[a21][b595][m595];
        end
    endgenerate
    generate 
        localparam integer b596 = 8;
        for (m596 = 0; m596 < 16; m596 = m596 + 1) 
        begin: inbit596
            assign data_11[m596 + b596*16 + a21*28*16] = data_11_array[a21][b596][m596];
        end
    endgenerate
    generate 
        localparam integer b597 = 9;
        for (m597 = 0; m597 < 16; m597 = m597 + 1) 
        begin: inbit597
            assign data_11[m597 + b597*16 + a21*28*16] = data_11_array[a21][b597][m597];
        end
    endgenerate
    generate 
        localparam integer b598 = 10;
        for (m598 = 0; m598 < 16; m598 = m598 + 1) 
        begin: inbit598
            assign data_11[m598 + b598*16 + a21*28*16] = data_11_array[a21][b598][m598];
        end
    endgenerate
    generate 
        localparam integer b599 = 11;
        for (m599 = 0; m599 < 16; m599 = m599 + 1) 
        begin: inbit599
            assign data_11[m599 + b599*16 + a21*28*16] = data_11_array[a21][b599][m599];
        end
    endgenerate
    generate 
        localparam integer b600 = 12;
        for (m600 = 0; m600 < 16; m600 = m600 + 1) 
        begin: inbit600
            assign data_11[m600 + b600*16 + a21*28*16] = data_11_array[a21][b600][m600];
        end
    endgenerate
    generate 
        localparam integer b601 = 13;
        for (m601 = 0; m601 < 16; m601 = m601 + 1) 
        begin: inbit601
            assign data_11[m601 + b601*16 + a21*28*16] = data_11_array[a21][b601][m601];
        end
    endgenerate
    generate 
        localparam integer b602 = 14;
        for (m602 = 0; m602 < 16; m602 = m602 + 1) 
        begin: inbit602
            assign data_11[m602 + b602*16 + a21*28*16] = data_11_array[a21][b602][m602];
        end
    endgenerate
    generate 
        localparam integer b603 = 15;
        for (m603 = 0; m603 < 16; m603 = m603 + 1) 
        begin: inbit603
            assign data_11[m603 + b603*16 + a21*28*16] = data_11_array[a21][b603][m603];
        end
    endgenerate
    generate 
        localparam integer b604 = 16;
        for (m604 = 0; m604 < 16; m604 = m604 + 1) 
        begin: inbit604
            assign data_11[m604 + b604*16 + a21*28*16] = data_11_array[a21][b604][m604];
        end
    endgenerate
    generate 
        localparam integer b605 = 17;
        for (m605 = 0; m605 < 16; m605 = m605 + 1) 
        begin: inbit605
            assign data_11[m605 + b605*16 + a21*28*16] = data_11_array[a21][b605][m605];
        end
    endgenerate
    generate 
        localparam integer b606 = 18;
        for (m606 = 0; m606 < 16; m606 = m606 + 1) 
        begin: inbit606
            assign data_11[m606 + b606*16 + a21*28*16] = data_11_array[a21][b606][m606];
        end
    endgenerate
    generate 
        localparam integer b607 = 19;
        for (m607 = 0; m607 < 16; m607 = m607 + 1) 
        begin: inbit607
            assign data_11[m607 + b607*16 + a21*28*16] = data_11_array[a21][b607][m607];
        end
    endgenerate
    generate 
        localparam integer b608 = 20;
        for (m608 = 0; m608 < 16; m608 = m608 + 1) 
        begin: inbit608
            assign data_11[m608 + b608*16 + a21*28*16] = data_11_array[a21][b608][m608];
        end
    endgenerate
    generate 
        localparam integer b609 = 21;
        for (m609 = 0; m609 < 16; m609 = m609 + 1) 
        begin: inbit609
            assign data_11[m609 + b609*16 + a21*28*16] = data_11_array[a21][b609][m609];
        end
    endgenerate
    generate 
        localparam integer b610 = 22;
        for (m610 = 0; m610 < 16; m610 = m610 + 1) 
        begin: inbit610
            assign data_11[m610 + b610*16 + a21*28*16] = data_11_array[a21][b610][m610];
        end
    endgenerate
    generate 
        localparam integer b611 = 23;
        for (m611 = 0; m611 < 16; m611 = m611 + 1) 
        begin: inbit611
            assign data_11[m611 + b611*16 + a21*28*16] = data_11_array[a21][b611][m611];
        end
    endgenerate
    generate 
        localparam integer b612 = 24;
        for (m612 = 0; m612 < 16; m612 = m612 + 1) 
        begin: inbit612
            assign data_11[m612 + b612*16 + a21*28*16] = data_11_array[a21][b612][m612];
        end
    endgenerate
    generate 
        localparam integer b613 = 25;
        for (m613 = 0; m613 < 16; m613 = m613 + 1) 
        begin: inbit613
            assign data_11[m613 + b613*16 + a21*28*16] = data_11_array[a21][b613][m613];
        end
    endgenerate
    generate 
        localparam integer b614 = 26;
        for (m614 = 0; m614 < 16; m614 = m614 + 1) 
        begin: inbit614
            assign data_11[m614 + b614*16 + a21*28*16] = data_11_array[a21][b614][m614];
        end
    endgenerate
    generate 
        localparam integer b615 = 27;
        for (m615 = 0; m615 < 16; m615 = m615 + 1) 
        begin: inbit615
            assign data_11[m615 + b615*16 + a21*28*16] = data_11_array[a21][b615][m615];
        end
    endgenerate
    localparam integer a22 = 22;
    generate 
        localparam integer b616 = 0;
        for (m616 = 0; m616 < 16; m616 = m616 + 1) 
        begin: inbit616
            assign data_11[m616 + b616*16 + a22*28*16] = data_11_array[a22][b616][m616];
        end
    endgenerate
    generate 
        localparam integer b617 = 1;
        for (m617 = 0; m617 < 16; m617 = m617 + 1) 
        begin: inbit617
            assign data_11[m617 + b617*16 + a22*28*16] = data_11_array[a22][b617][m617];
        end
    endgenerate
    generate 
        localparam integer b618 = 2;
        for (m618 = 0; m618 < 16; m618 = m618 + 1) 
        begin: inbit618
            assign data_11[m618 + b618*16 + a22*28*16] = data_11_array[a22][b618][m618];
        end
    endgenerate
    generate 
        localparam integer b619 = 3;
        for (m619 = 0; m619 < 16; m619 = m619 + 1) 
        begin: inbit619
            assign data_11[m619 + b619*16 + a22*28*16] = data_11_array[a22][b619][m619];
        end
    endgenerate
    generate 
        localparam integer b620 = 4;
        for (m620 = 0; m620 < 16; m620 = m620 + 1) 
        begin: inbit620
            assign data_11[m620 + b620*16 + a22*28*16] = data_11_array[a22][b620][m620];
        end
    endgenerate
    generate 
        localparam integer b621 = 5;
        for (m621 = 0; m621 < 16; m621 = m621 + 1) 
        begin: inbit621
            assign data_11[m621 + b621*16 + a22*28*16] = data_11_array[a22][b621][m621];
        end
    endgenerate
    generate 
        localparam integer b622 = 6;
        for (m622 = 0; m622 < 16; m622 = m622 + 1) 
        begin: inbit622
            assign data_11[m622 + b622*16 + a22*28*16] = data_11_array[a22][b622][m622];
        end
    endgenerate
    generate 
        localparam integer b623 = 7;
        for (m623 = 0; m623 < 16; m623 = m623 + 1) 
        begin: inbit623
            assign data_11[m623 + b623*16 + a22*28*16] = data_11_array[a22][b623][m623];
        end
    endgenerate
    generate 
        localparam integer b624 = 8;
        for (m624 = 0; m624 < 16; m624 = m624 + 1) 
        begin: inbit624
            assign data_11[m624 + b624*16 + a22*28*16] = data_11_array[a22][b624][m624];
        end
    endgenerate
    generate 
        localparam integer b625 = 9;
        for (m625 = 0; m625 < 16; m625 = m625 + 1) 
        begin: inbit625
            assign data_11[m625 + b625*16 + a22*28*16] = data_11_array[a22][b625][m625];
        end
    endgenerate
    generate 
        localparam integer b626 = 10;
        for (m626 = 0; m626 < 16; m626 = m626 + 1) 
        begin: inbit626
            assign data_11[m626 + b626*16 + a22*28*16] = data_11_array[a22][b626][m626];
        end
    endgenerate
    generate 
        localparam integer b627 = 11;
        for (m627 = 0; m627 < 16; m627 = m627 + 1) 
        begin: inbit627
            assign data_11[m627 + b627*16 + a22*28*16] = data_11_array[a22][b627][m627];
        end
    endgenerate
    generate 
        localparam integer b628 = 12;
        for (m628 = 0; m628 < 16; m628 = m628 + 1) 
        begin: inbit628
            assign data_11[m628 + b628*16 + a22*28*16] = data_11_array[a22][b628][m628];
        end
    endgenerate
    generate 
        localparam integer b629 = 13;
        for (m629 = 0; m629 < 16; m629 = m629 + 1) 
        begin: inbit629
            assign data_11[m629 + b629*16 + a22*28*16] = data_11_array[a22][b629][m629];
        end
    endgenerate
    generate 
        localparam integer b630 = 14;
        for (m630 = 0; m630 < 16; m630 = m630 + 1) 
        begin: inbit630
            assign data_11[m630 + b630*16 + a22*28*16] = data_11_array[a22][b630][m630];
        end
    endgenerate
    generate 
        localparam integer b631 = 15;
        for (m631 = 0; m631 < 16; m631 = m631 + 1) 
        begin: inbit631
            assign data_11[m631 + b631*16 + a22*28*16] = data_11_array[a22][b631][m631];
        end
    endgenerate
    generate 
        localparam integer b632 = 16;
        for (m632 = 0; m632 < 16; m632 = m632 + 1) 
        begin: inbit632
            assign data_11[m632 + b632*16 + a22*28*16] = data_11_array[a22][b632][m632];
        end
    endgenerate
    generate 
        localparam integer b633 = 17;
        for (m633 = 0; m633 < 16; m633 = m633 + 1) 
        begin: inbit633
            assign data_11[m633 + b633*16 + a22*28*16] = data_11_array[a22][b633][m633];
        end
    endgenerate
    generate 
        localparam integer b634 = 18;
        for (m634 = 0; m634 < 16; m634 = m634 + 1) 
        begin: inbit634
            assign data_11[m634 + b634*16 + a22*28*16] = data_11_array[a22][b634][m634];
        end
    endgenerate
    generate 
        localparam integer b635 = 19;
        for (m635 = 0; m635 < 16; m635 = m635 + 1) 
        begin: inbit635
            assign data_11[m635 + b635*16 + a22*28*16] = data_11_array[a22][b635][m635];
        end
    endgenerate
    generate 
        localparam integer b636 = 20;
        for (m636 = 0; m636 < 16; m636 = m636 + 1) 
        begin: inbit636
            assign data_11[m636 + b636*16 + a22*28*16] = data_11_array[a22][b636][m636];
        end
    endgenerate
    generate 
        localparam integer b637 = 21;
        for (m637 = 0; m637 < 16; m637 = m637 + 1) 
        begin: inbit637
            assign data_11[m637 + b637*16 + a22*28*16] = data_11_array[a22][b637][m637];
        end
    endgenerate
    generate 
        localparam integer b638 = 22;
        for (m638 = 0; m638 < 16; m638 = m638 + 1) 
        begin: inbit638
            assign data_11[m638 + b638*16 + a22*28*16] = data_11_array[a22][b638][m638];
        end
    endgenerate
    generate 
        localparam integer b639 = 23;
        for (m639 = 0; m639 < 16; m639 = m639 + 1) 
        begin: inbit639
            assign data_11[m639 + b639*16 + a22*28*16] = data_11_array[a22][b639][m639];
        end
    endgenerate
    generate 
        localparam integer b640 = 24;
        for (m640 = 0; m640 < 16; m640 = m640 + 1) 
        begin: inbit640
            assign data_11[m640 + b640*16 + a22*28*16] = data_11_array[a22][b640][m640];
        end
    endgenerate
    generate 
        localparam integer b641 = 25;
        for (m641 = 0; m641 < 16; m641 = m641 + 1) 
        begin: inbit641
            assign data_11[m641 + b641*16 + a22*28*16] = data_11_array[a22][b641][m641];
        end
    endgenerate
    generate 
        localparam integer b642 = 26;
        for (m642 = 0; m642 < 16; m642 = m642 + 1) 
        begin: inbit642
            assign data_11[m642 + b642*16 + a22*28*16] = data_11_array[a22][b642][m642];
        end
    endgenerate
    generate 
        localparam integer b643 = 27;
        for (m643 = 0; m643 < 16; m643 = m643 + 1) 
        begin: inbit643
            assign data_11[m643 + b643*16 + a22*28*16] = data_11_array[a22][b643][m643];
        end
    endgenerate
    localparam integer a23 = 23;
    generate 
        localparam integer b644 = 0;
        for (m644 = 0; m644 < 16; m644 = m644 + 1) 
        begin: inbit644
            assign data_11[m644 + b644*16 + a23*28*16] = data_11_array[a23][b644][m644];
        end
    endgenerate
    generate 
        localparam integer b645 = 1;
        for (m645 = 0; m645 < 16; m645 = m645 + 1) 
        begin: inbit645
            assign data_11[m645 + b645*16 + a23*28*16] = data_11_array[a23][b645][m645];
        end
    endgenerate
    generate 
        localparam integer b646 = 2;
        for (m646 = 0; m646 < 16; m646 = m646 + 1) 
        begin: inbit646
            assign data_11[m646 + b646*16 + a23*28*16] = data_11_array[a23][b646][m646];
        end
    endgenerate
    generate 
        localparam integer b647 = 3;
        for (m647 = 0; m647 < 16; m647 = m647 + 1) 
        begin: inbit647
            assign data_11[m647 + b647*16 + a23*28*16] = data_11_array[a23][b647][m647];
        end
    endgenerate
    generate 
        localparam integer b648 = 4;
        for (m648 = 0; m648 < 16; m648 = m648 + 1) 
        begin: inbit648
            assign data_11[m648 + b648*16 + a23*28*16] = data_11_array[a23][b648][m648];
        end
    endgenerate
    generate 
        localparam integer b649 = 5;
        for (m649 = 0; m649 < 16; m649 = m649 + 1) 
        begin: inbit649
            assign data_11[m649 + b649*16 + a23*28*16] = data_11_array[a23][b649][m649];
        end
    endgenerate
    generate 
        localparam integer b650 = 6;
        for (m650 = 0; m650 < 16; m650 = m650 + 1) 
        begin: inbit650
            assign data_11[m650 + b650*16 + a23*28*16] = data_11_array[a23][b650][m650];
        end
    endgenerate
    generate 
        localparam integer b651 = 7;
        for (m651 = 0; m651 < 16; m651 = m651 + 1) 
        begin: inbit651
            assign data_11[m651 + b651*16 + a23*28*16] = data_11_array[a23][b651][m651];
        end
    endgenerate
    generate 
        localparam integer b652 = 8;
        for (m652 = 0; m652 < 16; m652 = m652 + 1) 
        begin: inbit652
            assign data_11[m652 + b652*16 + a23*28*16] = data_11_array[a23][b652][m652];
        end
    endgenerate
    generate 
        localparam integer b653 = 9;
        for (m653 = 0; m653 < 16; m653 = m653 + 1) 
        begin: inbit653
            assign data_11[m653 + b653*16 + a23*28*16] = data_11_array[a23][b653][m653];
        end
    endgenerate
    generate 
        localparam integer b654 = 10;
        for (m654 = 0; m654 < 16; m654 = m654 + 1) 
        begin: inbit654
            assign data_11[m654 + b654*16 + a23*28*16] = data_11_array[a23][b654][m654];
        end
    endgenerate
    generate 
        localparam integer b655 = 11;
        for (m655 = 0; m655 < 16; m655 = m655 + 1) 
        begin: inbit655
            assign data_11[m655 + b655*16 + a23*28*16] = data_11_array[a23][b655][m655];
        end
    endgenerate
    generate 
        localparam integer b656 = 12;
        for (m656 = 0; m656 < 16; m656 = m656 + 1) 
        begin: inbit656
            assign data_11[m656 + b656*16 + a23*28*16] = data_11_array[a23][b656][m656];
        end
    endgenerate
    generate 
        localparam integer b657 = 13;
        for (m657 = 0; m657 < 16; m657 = m657 + 1) 
        begin: inbit657
            assign data_11[m657 + b657*16 + a23*28*16] = data_11_array[a23][b657][m657];
        end
    endgenerate
    generate 
        localparam integer b658 = 14;
        for (m658 = 0; m658 < 16; m658 = m658 + 1) 
        begin: inbit658
            assign data_11[m658 + b658*16 + a23*28*16] = data_11_array[a23][b658][m658];
        end
    endgenerate
    generate 
        localparam integer b659 = 15;
        for (m659 = 0; m659 < 16; m659 = m659 + 1) 
        begin: inbit659
            assign data_11[m659 + b659*16 + a23*28*16] = data_11_array[a23][b659][m659];
        end
    endgenerate
    generate 
        localparam integer b660 = 16;
        for (m660 = 0; m660 < 16; m660 = m660 + 1) 
        begin: inbit660
            assign data_11[m660 + b660*16 + a23*28*16] = data_11_array[a23][b660][m660];
        end
    endgenerate
    generate 
        localparam integer b661 = 17;
        for (m661 = 0; m661 < 16; m661 = m661 + 1) 
        begin: inbit661
            assign data_11[m661 + b661*16 + a23*28*16] = data_11_array[a23][b661][m661];
        end
    endgenerate
    generate 
        localparam integer b662 = 18;
        for (m662 = 0; m662 < 16; m662 = m662 + 1) 
        begin: inbit662
            assign data_11[m662 + b662*16 + a23*28*16] = data_11_array[a23][b662][m662];
        end
    endgenerate
    generate 
        localparam integer b663 = 19;
        for (m663 = 0; m663 < 16; m663 = m663 + 1) 
        begin: inbit663
            assign data_11[m663 + b663*16 + a23*28*16] = data_11_array[a23][b663][m663];
        end
    endgenerate
    generate 
        localparam integer b664 = 20;
        for (m664 = 0; m664 < 16; m664 = m664 + 1) 
        begin: inbit664
            assign data_11[m664 + b664*16 + a23*28*16] = data_11_array[a23][b664][m664];
        end
    endgenerate
    generate 
        localparam integer b665 = 21;
        for (m665 = 0; m665 < 16; m665 = m665 + 1) 
        begin: inbit665
            assign data_11[m665 + b665*16 + a23*28*16] = data_11_array[a23][b665][m665];
        end
    endgenerate
    generate 
        localparam integer b666 = 22;
        for (m666 = 0; m666 < 16; m666 = m666 + 1) 
        begin: inbit666
            assign data_11[m666 + b666*16 + a23*28*16] = data_11_array[a23][b666][m666];
        end
    endgenerate
    generate 
        localparam integer b667 = 23;
        for (m667 = 0; m667 < 16; m667 = m667 + 1) 
        begin: inbit667
            assign data_11[m667 + b667*16 + a23*28*16] = data_11_array[a23][b667][m667];
        end
    endgenerate
    generate 
        localparam integer b668 = 24;
        for (m668 = 0; m668 < 16; m668 = m668 + 1) 
        begin: inbit668
            assign data_11[m668 + b668*16 + a23*28*16] = data_11_array[a23][b668][m668];
        end
    endgenerate
    generate 
        localparam integer b669 = 25;
        for (m669 = 0; m669 < 16; m669 = m669 + 1) 
        begin: inbit669
            assign data_11[m669 + b669*16 + a23*28*16] = data_11_array[a23][b669][m669];
        end
    endgenerate
    generate 
        localparam integer b670 = 26;
        for (m670 = 0; m670 < 16; m670 = m670 + 1) 
        begin: inbit670
            assign data_11[m670 + b670*16 + a23*28*16] = data_11_array[a23][b670][m670];
        end
    endgenerate
    generate 
        localparam integer b671 = 27;
        for (m671 = 0; m671 < 16; m671 = m671 + 1) 
        begin: inbit671
            assign data_11[m671 + b671*16 + a23*28*16] = data_11_array[a23][b671][m671];
        end
    endgenerate
    localparam integer a24 = 24;
    generate 
        localparam integer b672 = 0;
        for (m672 = 0; m672 < 16; m672 = m672 + 1) 
        begin: inbit672
            assign data_11[m672 + b672*16 + a24*28*16] = data_11_array[a24][b672][m672];
        end
    endgenerate
    generate 
        localparam integer b673 = 1;
        for (m673 = 0; m673 < 16; m673 = m673 + 1) 
        begin: inbit673
            assign data_11[m673 + b673*16 + a24*28*16] = data_11_array[a24][b673][m673];
        end
    endgenerate
    generate 
        localparam integer b674 = 2;
        for (m674 = 0; m674 < 16; m674 = m674 + 1) 
        begin: inbit674
            assign data_11[m674 + b674*16 + a24*28*16] = data_11_array[a24][b674][m674];
        end
    endgenerate
    generate 
        localparam integer b675 = 3;
        for (m675 = 0; m675 < 16; m675 = m675 + 1) 
        begin: inbit675
            assign data_11[m675 + b675*16 + a24*28*16] = data_11_array[a24][b675][m675];
        end
    endgenerate
    generate 
        localparam integer b676 = 4;
        for (m676 = 0; m676 < 16; m676 = m676 + 1) 
        begin: inbit676
            assign data_11[m676 + b676*16 + a24*28*16] = data_11_array[a24][b676][m676];
        end
    endgenerate
    generate 
        localparam integer b677 = 5;
        for (m677 = 0; m677 < 16; m677 = m677 + 1) 
        begin: inbit677
            assign data_11[m677 + b677*16 + a24*28*16] = data_11_array[a24][b677][m677];
        end
    endgenerate
    generate 
        localparam integer b678 = 6;
        for (m678 = 0; m678 < 16; m678 = m678 + 1) 
        begin: inbit678
            assign data_11[m678 + b678*16 + a24*28*16] = data_11_array[a24][b678][m678];
        end
    endgenerate
    generate 
        localparam integer b679 = 7;
        for (m679 = 0; m679 < 16; m679 = m679 + 1) 
        begin: inbit679
            assign data_11[m679 + b679*16 + a24*28*16] = data_11_array[a24][b679][m679];
        end
    endgenerate
    generate 
        localparam integer b680 = 8;
        for (m680 = 0; m680 < 16; m680 = m680 + 1) 
        begin: inbit680
            assign data_11[m680 + b680*16 + a24*28*16] = data_11_array[a24][b680][m680];
        end
    endgenerate
    generate 
        localparam integer b681 = 9;
        for (m681 = 0; m681 < 16; m681 = m681 + 1) 
        begin: inbit681
            assign data_11[m681 + b681*16 + a24*28*16] = data_11_array[a24][b681][m681];
        end
    endgenerate
    generate 
        localparam integer b682 = 10;
        for (m682 = 0; m682 < 16; m682 = m682 + 1) 
        begin: inbit682
            assign data_11[m682 + b682*16 + a24*28*16] = data_11_array[a24][b682][m682];
        end
    endgenerate
    generate 
        localparam integer b683 = 11;
        for (m683 = 0; m683 < 16; m683 = m683 + 1) 
        begin: inbit683
            assign data_11[m683 + b683*16 + a24*28*16] = data_11_array[a24][b683][m683];
        end
    endgenerate
    generate 
        localparam integer b684 = 12;
        for (m684 = 0; m684 < 16; m684 = m684 + 1) 
        begin: inbit684
            assign data_11[m684 + b684*16 + a24*28*16] = data_11_array[a24][b684][m684];
        end
    endgenerate
    generate 
        localparam integer b685 = 13;
        for (m685 = 0; m685 < 16; m685 = m685 + 1) 
        begin: inbit685
            assign data_11[m685 + b685*16 + a24*28*16] = data_11_array[a24][b685][m685];
        end
    endgenerate
    generate 
        localparam integer b686 = 14;
        for (m686 = 0; m686 < 16; m686 = m686 + 1) 
        begin: inbit686
            assign data_11[m686 + b686*16 + a24*28*16] = data_11_array[a24][b686][m686];
        end
    endgenerate
    generate 
        localparam integer b687 = 15;
        for (m687 = 0; m687 < 16; m687 = m687 + 1) 
        begin: inbit687
            assign data_11[m687 + b687*16 + a24*28*16] = data_11_array[a24][b687][m687];
        end
    endgenerate
    generate 
        localparam integer b688 = 16;
        for (m688 = 0; m688 < 16; m688 = m688 + 1) 
        begin: inbit688
            assign data_11[m688 + b688*16 + a24*28*16] = data_11_array[a24][b688][m688];
        end
    endgenerate
    generate 
        localparam integer b689 = 17;
        for (m689 = 0; m689 < 16; m689 = m689 + 1) 
        begin: inbit689
            assign data_11[m689 + b689*16 + a24*28*16] = data_11_array[a24][b689][m689];
        end
    endgenerate
    generate 
        localparam integer b690 = 18;
        for (m690 = 0; m690 < 16; m690 = m690 + 1) 
        begin: inbit690
            assign data_11[m690 + b690*16 + a24*28*16] = data_11_array[a24][b690][m690];
        end
    endgenerate
    generate 
        localparam integer b691 = 19;
        for (m691 = 0; m691 < 16; m691 = m691 + 1) 
        begin: inbit691
            assign data_11[m691 + b691*16 + a24*28*16] = data_11_array[a24][b691][m691];
        end
    endgenerate
    generate 
        localparam integer b692 = 20;
        for (m692 = 0; m692 < 16; m692 = m692 + 1) 
        begin: inbit692
            assign data_11[m692 + b692*16 + a24*28*16] = data_11_array[a24][b692][m692];
        end
    endgenerate
    generate 
        localparam integer b693 = 21;
        for (m693 = 0; m693 < 16; m693 = m693 + 1) 
        begin: inbit693
            assign data_11[m693 + b693*16 + a24*28*16] = data_11_array[a24][b693][m693];
        end
    endgenerate
    generate 
        localparam integer b694 = 22;
        for (m694 = 0; m694 < 16; m694 = m694 + 1) 
        begin: inbit694
            assign data_11[m694 + b694*16 + a24*28*16] = data_11_array[a24][b694][m694];
        end
    endgenerate
    generate 
        localparam integer b695 = 23;
        for (m695 = 0; m695 < 16; m695 = m695 + 1) 
        begin: inbit695
            assign data_11[m695 + b695*16 + a24*28*16] = data_11_array[a24][b695][m695];
        end
    endgenerate
    generate 
        localparam integer b696 = 24;
        for (m696 = 0; m696 < 16; m696 = m696 + 1) 
        begin: inbit696
            assign data_11[m696 + b696*16 + a24*28*16] = data_11_array[a24][b696][m696];
        end
    endgenerate
    generate 
        localparam integer b697 = 25;
        for (m697 = 0; m697 < 16; m697 = m697 + 1) 
        begin: inbit697
            assign data_11[m697 + b697*16 + a24*28*16] = data_11_array[a24][b697][m697];
        end
    endgenerate
    generate 
        localparam integer b698 = 26;
        for (m698 = 0; m698 < 16; m698 = m698 + 1) 
        begin: inbit698
            assign data_11[m698 + b698*16 + a24*28*16] = data_11_array[a24][b698][m698];
        end
    endgenerate
    generate 
        localparam integer b699 = 27;
        for (m699 = 0; m699 < 16; m699 = m699 + 1) 
        begin: inbit699
            assign data_11[m699 + b699*16 + a24*28*16] = data_11_array[a24][b699][m699];
        end
    endgenerate
    localparam integer a25 = 25;
    generate 
        localparam integer b700 = 0;
        for (m700 = 0; m700 < 16; m700 = m700 + 1) 
        begin: inbit700
            assign data_11[m700 + b700*16 + a25*28*16] = data_11_array[a25][b700][m700];
        end
    endgenerate
    generate 
        localparam integer b701 = 1;
        for (m701 = 0; m701 < 16; m701 = m701 + 1) 
        begin: inbit701
            assign data_11[m701 + b701*16 + a25*28*16] = data_11_array[a25][b701][m701];
        end
    endgenerate
    generate 
        localparam integer b702 = 2;
        for (m702 = 0; m702 < 16; m702 = m702 + 1) 
        begin: inbit702
            assign data_11[m702 + b702*16 + a25*28*16] = data_11_array[a25][b702][m702];
        end
    endgenerate
    generate 
        localparam integer b703 = 3;
        for (m703 = 0; m703 < 16; m703 = m703 + 1) 
        begin: inbit703
            assign data_11[m703 + b703*16 + a25*28*16] = data_11_array[a25][b703][m703];
        end
    endgenerate
    generate 
        localparam integer b704 = 4;
        for (m704 = 0; m704 < 16; m704 = m704 + 1) 
        begin: inbit704
            assign data_11[m704 + b704*16 + a25*28*16] = data_11_array[a25][b704][m704];
        end
    endgenerate
    generate 
        localparam integer b705 = 5;
        for (m705 = 0; m705 < 16; m705 = m705 + 1) 
        begin: inbit705
            assign data_11[m705 + b705*16 + a25*28*16] = data_11_array[a25][b705][m705];
        end
    endgenerate
    generate 
        localparam integer b706 = 6;
        for (m706 = 0; m706 < 16; m706 = m706 + 1) 
        begin: inbit706
            assign data_11[m706 + b706*16 + a25*28*16] = data_11_array[a25][b706][m706];
        end
    endgenerate
    generate 
        localparam integer b707 = 7;
        for (m707 = 0; m707 < 16; m707 = m707 + 1) 
        begin: inbit707
            assign data_11[m707 + b707*16 + a25*28*16] = data_11_array[a25][b707][m707];
        end
    endgenerate
    generate 
        localparam integer b708 = 8;
        for (m708 = 0; m708 < 16; m708 = m708 + 1) 
        begin: inbit708
            assign data_11[m708 + b708*16 + a25*28*16] = data_11_array[a25][b708][m708];
        end
    endgenerate
    generate 
        localparam integer b709 = 9;
        for (m709 = 0; m709 < 16; m709 = m709 + 1) 
        begin: inbit709
            assign data_11[m709 + b709*16 + a25*28*16] = data_11_array[a25][b709][m709];
        end
    endgenerate
    generate 
        localparam integer b710 = 10;
        for (m710 = 0; m710 < 16; m710 = m710 + 1) 
        begin: inbit710
            assign data_11[m710 + b710*16 + a25*28*16] = data_11_array[a25][b710][m710];
        end
    endgenerate
    generate 
        localparam integer b711 = 11;
        for (m711 = 0; m711 < 16; m711 = m711 + 1) 
        begin: inbit711
            assign data_11[m711 + b711*16 + a25*28*16] = data_11_array[a25][b711][m711];
        end
    endgenerate
    generate 
        localparam integer b712 = 12;
        for (m712 = 0; m712 < 16; m712 = m712 + 1) 
        begin: inbit712
            assign data_11[m712 + b712*16 + a25*28*16] = data_11_array[a25][b712][m712];
        end
    endgenerate
    generate 
        localparam integer b713 = 13;
        for (m713 = 0; m713 < 16; m713 = m713 + 1) 
        begin: inbit713
            assign data_11[m713 + b713*16 + a25*28*16] = data_11_array[a25][b713][m713];
        end
    endgenerate
    generate 
        localparam integer b714 = 14;
        for (m714 = 0; m714 < 16; m714 = m714 + 1) 
        begin: inbit714
            assign data_11[m714 + b714*16 + a25*28*16] = data_11_array[a25][b714][m714];
        end
    endgenerate
    generate 
        localparam integer b715 = 15;
        for (m715 = 0; m715 < 16; m715 = m715 + 1) 
        begin: inbit715
            assign data_11[m715 + b715*16 + a25*28*16] = data_11_array[a25][b715][m715];
        end
    endgenerate
    generate 
        localparam integer b716 = 16;
        for (m716 = 0; m716 < 16; m716 = m716 + 1) 
        begin: inbit716
            assign data_11[m716 + b716*16 + a25*28*16] = data_11_array[a25][b716][m716];
        end
    endgenerate
    generate 
        localparam integer b717 = 17;
        for (m717 = 0; m717 < 16; m717 = m717 + 1) 
        begin: inbit717
            assign data_11[m717 + b717*16 + a25*28*16] = data_11_array[a25][b717][m717];
        end
    endgenerate
    generate 
        localparam integer b718 = 18;
        for (m718 = 0; m718 < 16; m718 = m718 + 1) 
        begin: inbit718
            assign data_11[m718 + b718*16 + a25*28*16] = data_11_array[a25][b718][m718];
        end
    endgenerate
    generate 
        localparam integer b719 = 19;
        for (m719 = 0; m719 < 16; m719 = m719 + 1) 
        begin: inbit719
            assign data_11[m719 + b719*16 + a25*28*16] = data_11_array[a25][b719][m719];
        end
    endgenerate
    generate 
        localparam integer b720 = 20;
        for (m720 = 0; m720 < 16; m720 = m720 + 1) 
        begin: inbit720
            assign data_11[m720 + b720*16 + a25*28*16] = data_11_array[a25][b720][m720];
        end
    endgenerate
    generate 
        localparam integer b721 = 21;
        for (m721 = 0; m721 < 16; m721 = m721 + 1) 
        begin: inbit721
            assign data_11[m721 + b721*16 + a25*28*16] = data_11_array[a25][b721][m721];
        end
    endgenerate
    generate 
        localparam integer b722 = 22;
        for (m722 = 0; m722 < 16; m722 = m722 + 1) 
        begin: inbit722
            assign data_11[m722 + b722*16 + a25*28*16] = data_11_array[a25][b722][m722];
        end
    endgenerate
    generate 
        localparam integer b723 = 23;
        for (m723 = 0; m723 < 16; m723 = m723 + 1) 
        begin: inbit723
            assign data_11[m723 + b723*16 + a25*28*16] = data_11_array[a25][b723][m723];
        end
    endgenerate
    generate 
        localparam integer b724 = 24;
        for (m724 = 0; m724 < 16; m724 = m724 + 1) 
        begin: inbit724
            assign data_11[m724 + b724*16 + a25*28*16] = data_11_array[a25][b724][m724];
        end
    endgenerate
    generate 
        localparam integer b725 = 25;
        for (m725 = 0; m725 < 16; m725 = m725 + 1) 
        begin: inbit725
            assign data_11[m725 + b725*16 + a25*28*16] = data_11_array[a25][b725][m725];
        end
    endgenerate
    generate 
        localparam integer b726 = 26;
        for (m726 = 0; m726 < 16; m726 = m726 + 1) 
        begin: inbit726
            assign data_11[m726 + b726*16 + a25*28*16] = data_11_array[a25][b726][m726];
        end
    endgenerate
    generate 
        localparam integer b727 = 27;
        for (m727 = 0; m727 < 16; m727 = m727 + 1) 
        begin: inbit727
            assign data_11[m727 + b727*16 + a25*28*16] = data_11_array[a25][b727][m727];
        end
    endgenerate
    localparam integer a26 = 26;
    generate 
        localparam integer b728 = 0;
        for (m728 = 0; m728 < 16; m728 = m728 + 1) 
        begin: inbit728
            assign data_11[m728 + b728*16 + a26*28*16] = data_11_array[a26][b728][m728];
        end
    endgenerate
    generate 
        localparam integer b729 = 1;
        for (m729 = 0; m729 < 16; m729 = m729 + 1) 
        begin: inbit729
            assign data_11[m729 + b729*16 + a26*28*16] = data_11_array[a26][b729][m729];
        end
    endgenerate
    generate 
        localparam integer b730 = 2;
        for (m730 = 0; m730 < 16; m730 = m730 + 1) 
        begin: inbit730
            assign data_11[m730 + b730*16 + a26*28*16] = data_11_array[a26][b730][m730];
        end
    endgenerate
    generate 
        localparam integer b731 = 3;
        for (m731 = 0; m731 < 16; m731 = m731 + 1) 
        begin: inbit731
            assign data_11[m731 + b731*16 + a26*28*16] = data_11_array[a26][b731][m731];
        end
    endgenerate
    generate 
        localparam integer b732 = 4;
        for (m732 = 0; m732 < 16; m732 = m732 + 1) 
        begin: inbit732
            assign data_11[m732 + b732*16 + a26*28*16] = data_11_array[a26][b732][m732];
        end
    endgenerate
    generate 
        localparam integer b733 = 5;
        for (m733 = 0; m733 < 16; m733 = m733 + 1) 
        begin: inbit733
            assign data_11[m733 + b733*16 + a26*28*16] = data_11_array[a26][b733][m733];
        end
    endgenerate
    generate 
        localparam integer b734 = 6;
        for (m734 = 0; m734 < 16; m734 = m734 + 1) 
        begin: inbit734
            assign data_11[m734 + b734*16 + a26*28*16] = data_11_array[a26][b734][m734];
        end
    endgenerate
    generate 
        localparam integer b735 = 7;
        for (m735 = 0; m735 < 16; m735 = m735 + 1) 
        begin: inbit735
            assign data_11[m735 + b735*16 + a26*28*16] = data_11_array[a26][b735][m735];
        end
    endgenerate
    generate 
        localparam integer b736 = 8;
        for (m736 = 0; m736 < 16; m736 = m736 + 1) 
        begin: inbit736
            assign data_11[m736 + b736*16 + a26*28*16] = data_11_array[a26][b736][m736];
        end
    endgenerate
    generate 
        localparam integer b737 = 9;
        for (m737 = 0; m737 < 16; m737 = m737 + 1) 
        begin: inbit737
            assign data_11[m737 + b737*16 + a26*28*16] = data_11_array[a26][b737][m737];
        end
    endgenerate
    generate 
        localparam integer b738 = 10;
        for (m738 = 0; m738 < 16; m738 = m738 + 1) 
        begin: inbit738
            assign data_11[m738 + b738*16 + a26*28*16] = data_11_array[a26][b738][m738];
        end
    endgenerate
    generate 
        localparam integer b739 = 11;
        for (m739 = 0; m739 < 16; m739 = m739 + 1) 
        begin: inbit739
            assign data_11[m739 + b739*16 + a26*28*16] = data_11_array[a26][b739][m739];
        end
    endgenerate
    generate 
        localparam integer b740 = 12;
        for (m740 = 0; m740 < 16; m740 = m740 + 1) 
        begin: inbit740
            assign data_11[m740 + b740*16 + a26*28*16] = data_11_array[a26][b740][m740];
        end
    endgenerate
    generate 
        localparam integer b741 = 13;
        for (m741 = 0; m741 < 16; m741 = m741 + 1) 
        begin: inbit741
            assign data_11[m741 + b741*16 + a26*28*16] = data_11_array[a26][b741][m741];
        end
    endgenerate
    generate 
        localparam integer b742 = 14;
        for (m742 = 0; m742 < 16; m742 = m742 + 1) 
        begin: inbit742
            assign data_11[m742 + b742*16 + a26*28*16] = data_11_array[a26][b742][m742];
        end
    endgenerate
    generate 
        localparam integer b743 = 15;
        for (m743 = 0; m743 < 16; m743 = m743 + 1) 
        begin: inbit743
            assign data_11[m743 + b743*16 + a26*28*16] = data_11_array[a26][b743][m743];
        end
    endgenerate
    generate 
        localparam integer b744 = 16;
        for (m744 = 0; m744 < 16; m744 = m744 + 1) 
        begin: inbit744
            assign data_11[m744 + b744*16 + a26*28*16] = data_11_array[a26][b744][m744];
        end
    endgenerate
    generate 
        localparam integer b745 = 17;
        for (m745 = 0; m745 < 16; m745 = m745 + 1) 
        begin: inbit745
            assign data_11[m745 + b745*16 + a26*28*16] = data_11_array[a26][b745][m745];
        end
    endgenerate
    generate 
        localparam integer b746 = 18;
        for (m746 = 0; m746 < 16; m746 = m746 + 1) 
        begin: inbit746
            assign data_11[m746 + b746*16 + a26*28*16] = data_11_array[a26][b746][m746];
        end
    endgenerate
    generate 
        localparam integer b747 = 19;
        for (m747 = 0; m747 < 16; m747 = m747 + 1) 
        begin: inbit747
            assign data_11[m747 + b747*16 + a26*28*16] = data_11_array[a26][b747][m747];
        end
    endgenerate
    generate 
        localparam integer b748 = 20;
        for (m748 = 0; m748 < 16; m748 = m748 + 1) 
        begin: inbit748
            assign data_11[m748 + b748*16 + a26*28*16] = data_11_array[a26][b748][m748];
        end
    endgenerate
    generate 
        localparam integer b749 = 21;
        for (m749 = 0; m749 < 16; m749 = m749 + 1) 
        begin: inbit749
            assign data_11[m749 + b749*16 + a26*28*16] = data_11_array[a26][b749][m749];
        end
    endgenerate
    generate 
        localparam integer b750 = 22;
        for (m750 = 0; m750 < 16; m750 = m750 + 1) 
        begin: inbit750
            assign data_11[m750 + b750*16 + a26*28*16] = data_11_array[a26][b750][m750];
        end
    endgenerate
    generate 
        localparam integer b751 = 23;
        for (m751 = 0; m751 < 16; m751 = m751 + 1) 
        begin: inbit751
            assign data_11[m751 + b751*16 + a26*28*16] = data_11_array[a26][b751][m751];
        end
    endgenerate
    generate 
        localparam integer b752 = 24;
        for (m752 = 0; m752 < 16; m752 = m752 + 1) 
        begin: inbit752
            assign data_11[m752 + b752*16 + a26*28*16] = data_11_array[a26][b752][m752];
        end
    endgenerate
    generate 
        localparam integer b753 = 25;
        for (m753 = 0; m753 < 16; m753 = m753 + 1) 
        begin: inbit753
            assign data_11[m753 + b753*16 + a26*28*16] = data_11_array[a26][b753][m753];
        end
    endgenerate
    generate 
        localparam integer b754 = 26;
        for (m754 = 0; m754 < 16; m754 = m754 + 1) 
        begin: inbit754
            assign data_11[m754 + b754*16 + a26*28*16] = data_11_array[a26][b754][m754];
        end
    endgenerate
    generate 
        localparam integer b755 = 27;
        for (m755 = 0; m755 < 16; m755 = m755 + 1) 
        begin: inbit755
            assign data_11[m755 + b755*16 + a26*28*16] = data_11_array[a26][b755][m755];
        end
    endgenerate
    localparam integer a27 = 27;
    generate 
        localparam integer b756 = 0;
        for (m756 = 0; m756 < 16; m756 = m756 + 1) 
        begin: inbit756
            assign data_11[m756 + b756*16 + a27*28*16] = data_11_array[a27][b756][m756];
        end
    endgenerate
    generate 
        localparam integer b757 = 1;
        for (m757 = 0; m757 < 16; m757 = m757 + 1) 
        begin: inbit757
            assign data_11[m757 + b757*16 + a27*28*16] = data_11_array[a27][b757][m757];
        end
    endgenerate
    generate 
        localparam integer b758 = 2;
        for (m758 = 0; m758 < 16; m758 = m758 + 1) 
        begin: inbit758
            assign data_11[m758 + b758*16 + a27*28*16] = data_11_array[a27][b758][m758];
        end
    endgenerate
    generate 
        localparam integer b759 = 3;
        for (m759 = 0; m759 < 16; m759 = m759 + 1) 
        begin: inbit759
            assign data_11[m759 + b759*16 + a27*28*16] = data_11_array[a27][b759][m759];
        end
    endgenerate
    generate 
        localparam integer b760 = 4;
        for (m760 = 0; m760 < 16; m760 = m760 + 1) 
        begin: inbit760
            assign data_11[m760 + b760*16 + a27*28*16] = data_11_array[a27][b760][m760];
        end
    endgenerate
    generate 
        localparam integer b761 = 5;
        for (m761 = 0; m761 < 16; m761 = m761 + 1) 
        begin: inbit761
            assign data_11[m761 + b761*16 + a27*28*16] = data_11_array[a27][b761][m761];
        end
    endgenerate
    generate 
        localparam integer b762 = 6;
        for (m762 = 0; m762 < 16; m762 = m762 + 1) 
        begin: inbit762
            assign data_11[m762 + b762*16 + a27*28*16] = data_11_array[a27][b762][m762];
        end
    endgenerate
    generate 
        localparam integer b763 = 7;
        for (m763 = 0; m763 < 16; m763 = m763 + 1) 
        begin: inbit763
            assign data_11[m763 + b763*16 + a27*28*16] = data_11_array[a27][b763][m763];
        end
    endgenerate
    generate 
        localparam integer b764 = 8;
        for (m764 = 0; m764 < 16; m764 = m764 + 1) 
        begin: inbit764
            assign data_11[m764 + b764*16 + a27*28*16] = data_11_array[a27][b764][m764];
        end
    endgenerate
    generate 
        localparam integer b765 = 9;
        for (m765 = 0; m765 < 16; m765 = m765 + 1) 
        begin: inbit765
            assign data_11[m765 + b765*16 + a27*28*16] = data_11_array[a27][b765][m765];
        end
    endgenerate
    generate 
        localparam integer b766 = 10;
        for (m766 = 0; m766 < 16; m766 = m766 + 1) 
        begin: inbit766
            assign data_11[m766 + b766*16 + a27*28*16] = data_11_array[a27][b766][m766];
        end
    endgenerate
    generate 
        localparam integer b767 = 11;
        for (m767 = 0; m767 < 16; m767 = m767 + 1) 
        begin: inbit767
            assign data_11[m767 + b767*16 + a27*28*16] = data_11_array[a27][b767][m767];
        end
    endgenerate
    generate 
        localparam integer b768 = 12;
        for (m768 = 0; m768 < 16; m768 = m768 + 1) 
        begin: inbit768
            assign data_11[m768 + b768*16 + a27*28*16] = data_11_array[a27][b768][m768];
        end
    endgenerate
    generate 
        localparam integer b769 = 13;
        for (m769 = 0; m769 < 16; m769 = m769 + 1) 
        begin: inbit769
            assign data_11[m769 + b769*16 + a27*28*16] = data_11_array[a27][b769][m769];
        end
    endgenerate
    generate 
        localparam integer b770 = 14;
        for (m770 = 0; m770 < 16; m770 = m770 + 1) 
        begin: inbit770
            assign data_11[m770 + b770*16 + a27*28*16] = data_11_array[a27][b770][m770];
        end
    endgenerate
    generate 
        localparam integer b771 = 15;
        for (m771 = 0; m771 < 16; m771 = m771 + 1) 
        begin: inbit771
            assign data_11[m771 + b771*16 + a27*28*16] = data_11_array[a27][b771][m771];
        end
    endgenerate
    generate 
        localparam integer b772 = 16;
        for (m772 = 0; m772 < 16; m772 = m772 + 1) 
        begin: inbit772
            assign data_11[m772 + b772*16 + a27*28*16] = data_11_array[a27][b772][m772];
        end
    endgenerate
    generate 
        localparam integer b773 = 17;
        for (m773 = 0; m773 < 16; m773 = m773 + 1) 
        begin: inbit773
            assign data_11[m773 + b773*16 + a27*28*16] = data_11_array[a27][b773][m773];
        end
    endgenerate
    generate 
        localparam integer b774 = 18;
        for (m774 = 0; m774 < 16; m774 = m774 + 1) 
        begin: inbit774
            assign data_11[m774 + b774*16 + a27*28*16] = data_11_array[a27][b774][m774];
        end
    endgenerate
    generate 
        localparam integer b775 = 19;
        for (m775 = 0; m775 < 16; m775 = m775 + 1) 
        begin: inbit775
            assign data_11[m775 + b775*16 + a27*28*16] = data_11_array[a27][b775][m775];
        end
    endgenerate
    generate 
        localparam integer b776 = 20;
        for (m776 = 0; m776 < 16; m776 = m776 + 1) 
        begin: inbit776
            assign data_11[m776 + b776*16 + a27*28*16] = data_11_array[a27][b776][m776];
        end
    endgenerate
    generate 
        localparam integer b777 = 21;
        for (m777 = 0; m777 < 16; m777 = m777 + 1) 
        begin: inbit777
            assign data_11[m777 + b777*16 + a27*28*16] = data_11_array[a27][b777][m777];
        end
    endgenerate
    generate 
        localparam integer b778 = 22;
        for (m778 = 0; m778 < 16; m778 = m778 + 1) 
        begin: inbit778
            assign data_11[m778 + b778*16 + a27*28*16] = data_11_array[a27][b778][m778];
        end
    endgenerate
    generate 
        localparam integer b779 = 23;
        for (m779 = 0; m779 < 16; m779 = m779 + 1) 
        begin: inbit779
            assign data_11[m779 + b779*16 + a27*28*16] = data_11_array[a27][b779][m779];
        end
    endgenerate
    generate 
        localparam integer b780 = 24;
        for (m780 = 0; m780 < 16; m780 = m780 + 1) 
        begin: inbit780
            assign data_11[m780 + b780*16 + a27*28*16] = data_11_array[a27][b780][m780];
        end
    endgenerate
    generate 
        localparam integer b781 = 25;
        for (m781 = 0; m781 < 16; m781 = m781 + 1) 
        begin: inbit781
            assign data_11[m781 + b781*16 + a27*28*16] = data_11_array[a27][b781][m781];
        end
    endgenerate
    generate 
        localparam integer b782 = 26;
        for (m782 = 0; m782 < 16; m782 = m782 + 1) 
        begin: inbit782
            assign data_11[m782 + b782*16 + a27*28*16] = data_11_array[a27][b782][m782];
        end
    endgenerate
    generate 
        localparam integer b783 = 27;
        for (m783 = 0; m783 < 16; m783 = m783 + 1) 
        begin: inbit783
            assign data_11[m783 + b783*16 + a27*28*16] = data_11_array[a27][b783][m783];
        end
    endgenerate
  
  ////ROW 0
  generate
    localparam integer j0 = 0;
    for (i0 = 0; i0 < 24; i0 = i0 + 1)
    begin: addbit0
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j0+0][i0+0]), .Out(multi0[0][i0]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j0+0][i0+1]), .Out(multi0[1][i0]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j0+0][i0+2]), .Out(multi0[2][i0]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j0+0][i0+3]), .Out(multi0[3][i0]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j0+0][i0+4]), .Out(multi0[4][i0]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j0+1][i0+0]), .Out(multi0[5][i0]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j0+1][i0+1]), .Out(multi0[6][i0]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j0+1][i0+2]), .Out(multi0[7][i0]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j0+1][i0+3]), .Out(multi0[8][i0]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j0+1][i0+4]), .Out(multi0[9][i0]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j0+2][i0+0]), .Out(multi0[10][i0]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j0+2][i0+1]), .Out(multi0[11][i0]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j0+2][i0+2]), .Out(multi0[12][i0]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j0+2][i0+3]), .Out(multi0[13][i0]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j0+2][i0+4]), .Out(multi0[14][i0]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j0+3][i0+0]), .Out(multi0[15][i0]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j0+3][i0+1]), .Out(multi0[16][i0]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j0+3][i0+2]), .Out(multi0[17][i0]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j0+3][i0+3]), .Out(multi0[18][i0]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j0+3][i0+4]), .Out(multi0[19][i0]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j0+4][i0+0]), .Out(multi0[20][i0]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j0+4][i0+1]), .Out(multi0[21][i0]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j0+4][i0+2]), .Out(multi0[22][i0]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j0+4][i0+3]), .Out(multi0[23][i0]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j0+4][i0+4]), .Out(multi0[24][i0]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi0[0][i0]), .B(multi0[1][i0]), .Out(sum0[0][i0]));
      FP16_Add stage026(.A(multi0[2][i0]), .B(multi0[3][i0]), .Out(sum0[1][i0]));
      FP16_Add stage027(.A(multi0[4][i0]), .B(multi0[5][i0]), .Out(sum0[2][i0]));
      FP16_Add stage028(.A(multi0[6][i0]), .B(multi0[7][i0]), .Out(sum0[3][i0]));
      FP16_Add stage029(.A(multi0[8][i0]), .B(multi0[9][i0]), .Out(sum0[4][i0]));
      FP16_Add stage030(.A(multi0[10][i0]), .B(multi0[11][i0]), .Out(sum0[5][i0]));
      FP16_Add stage031(.A(multi0[12][i0]), .B(multi0[13][i0]), .Out(sum0[6][i0]));
      FP16_Add stage032(.A(multi0[14][i0]), .B(multi0[15][i0]), .Out(sum0[7][i0]));
      FP16_Add stage033(.A(multi0[16][i0]), .B(multi0[17][i0]), .Out(sum0[8][i0]));
      FP16_Add stage034(.A(multi0[18][i0]), .B(multi0[19][i0]), .Out(sum0[9][i0]));
      FP16_Add stage035(.A(multi0[20][i0]), .B(multi0[21][i0]), .Out(sum0[10][i0]));
      FP16_Add stage036(.A(multi0[22][i0]), .B(multi0[23][i0]), .Out(sum0[11][i0]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum0[0][i0]), .B(sum0[1][i0]), .Out(sum0[12][i0]));
      FP16_Add stage038(.A(sum0[2][i0]), .B(sum0[3][i0]), .Out(sum0[13][i0]));
      FP16_Add stage039(.A(sum0[4][i0]), .B(sum0[5][i0]), .Out(sum0[14][i0]));
      FP16_Add stage040(.A(sum0[6][i0]), .B(sum0[7][i0]), .Out(sum0[15][i0]));
      FP16_Add stage041(.A(sum0[8][i0]), .B(sum0[9][i0]), .Out(sum0[16][i0]));
      FP16_Add stage042(.A(sum0[10][i0]), .B(sum0[11][i0]), .Out(sum0[17][i0]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum0[12][i0]), .B(sum0[13][i0]), .Out(sum0[18][i0]));
      FP16_Add stage044(.A(sum0[14][i0]), .B(sum0[15][i0]), .Out(sum0[19][i0]));
      FP16_Add stage045(.A(sum0[16][i0]), .B(sum0[17][i0]), .Out(sum0[20][i0]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum0[18][i0]), .B(sum0[19][i0]), .Out(sum0[21][i0]));
      FP16_Add stage047(.A(sum0[20][i0]), .B(multi0[24][i0]), .Out(sum0[22][i0]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum0[21][i0]), .B(sum0[22][i0]), .Out(sum0[23][i0]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum0[23][i0]), .B(feature4Bias), .Out(data_11_array[j0][i0]));
    end
  endgenerate
  
  ////ROW 1
  generate
    localparam integer j1 = 1;
    for (i1 = 0; i1 < 24; i1 = i1 + 1)
    begin: addbit1
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j1+0][i1+0]), .Out(multi1[0][i1]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j1+0][i1+1]), .Out(multi1[1][i1]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j1+0][i1+2]), .Out(multi1[2][i1]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j1+0][i1+3]), .Out(multi1[3][i1]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j1+0][i1+4]), .Out(multi1[4][i1]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j1+1][i1+0]), .Out(multi1[5][i1]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j1+1][i1+1]), .Out(multi1[6][i1]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j1+1][i1+2]), .Out(multi1[7][i1]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j1+1][i1+3]), .Out(multi1[8][i1]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j1+1][i1+4]), .Out(multi1[9][i1]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j1+2][i1+0]), .Out(multi1[10][i1]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j1+2][i1+1]), .Out(multi1[11][i1]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j1+2][i1+2]), .Out(multi1[12][i1]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j1+2][i1+3]), .Out(multi1[13][i1]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j1+2][i1+4]), .Out(multi1[14][i1]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j1+3][i1+0]), .Out(multi1[15][i1]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j1+3][i1+1]), .Out(multi1[16][i1]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j1+3][i1+2]), .Out(multi1[17][i1]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j1+3][i1+3]), .Out(multi1[18][i1]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j1+3][i1+4]), .Out(multi1[19][i1]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j1+4][i1+0]), .Out(multi1[20][i1]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j1+4][i1+1]), .Out(multi1[21][i1]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j1+4][i1+2]), .Out(multi1[22][i1]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j1+4][i1+3]), .Out(multi1[23][i1]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j1+4][i1+4]), .Out(multi1[24][i1]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi1[0][i1]), .B(multi1[1][i1]), .Out(sum1[0][i1]));
      FP16_Add stage026(.A(multi1[2][i1]), .B(multi1[3][i1]), .Out(sum1[1][i1]));
      FP16_Add stage027(.A(multi1[4][i1]), .B(multi1[5][i1]), .Out(sum1[2][i1]));
      FP16_Add stage028(.A(multi1[6][i1]), .B(multi1[7][i1]), .Out(sum1[3][i1]));
      FP16_Add stage029(.A(multi1[8][i1]), .B(multi1[9][i1]), .Out(sum1[4][i1]));
      FP16_Add stage030(.A(multi1[10][i1]), .B(multi1[11][i1]), .Out(sum1[5][i1]));
      FP16_Add stage031(.A(multi1[12][i1]), .B(multi1[13][i1]), .Out(sum1[6][i1]));
      FP16_Add stage032(.A(multi1[14][i1]), .B(multi1[15][i1]), .Out(sum1[7][i1]));
      FP16_Add stage033(.A(multi1[16][i1]), .B(multi1[17][i1]), .Out(sum1[8][i1]));
      FP16_Add stage034(.A(multi1[18][i1]), .B(multi1[19][i1]), .Out(sum1[9][i1]));
      FP16_Add stage035(.A(multi1[20][i1]), .B(multi1[21][i1]), .Out(sum1[10][i1]));
      FP16_Add stage036(.A(multi1[22][i1]), .B(multi1[23][i1]), .Out(sum1[11][i1]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum1[0][i1]), .B(sum1[1][i1]), .Out(sum1[12][i1]));
      FP16_Add stage038(.A(sum1[2][i1]), .B(sum1[3][i1]), .Out(sum1[13][i1]));
      FP16_Add stage039(.A(sum1[4][i1]), .B(sum1[5][i1]), .Out(sum1[14][i1]));
      FP16_Add stage040(.A(sum1[6][i1]), .B(sum1[7][i1]), .Out(sum1[15][i1]));
      FP16_Add stage041(.A(sum1[8][i1]), .B(sum1[9][i1]), .Out(sum1[16][i1]));
      FP16_Add stage042(.A(sum1[10][i1]), .B(sum1[11][i1]), .Out(sum1[17][i1]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum1[12][i1]), .B(sum1[13][i1]), .Out(sum1[18][i1]));
      FP16_Add stage044(.A(sum1[14][i1]), .B(sum1[15][i1]), .Out(sum1[19][i1]));
      FP16_Add stage045(.A(sum1[16][i1]), .B(sum1[17][i1]), .Out(sum1[20][i1]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum1[18][i1]), .B(sum1[19][i1]), .Out(sum1[21][i1]));
      FP16_Add stage047(.A(sum1[20][i1]), .B(multi1[24][i1]), .Out(sum1[22][i1]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum1[21][i1]), .B(sum1[22][i1]), .Out(sum1[23][i1]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum1[23][i1]), .B(feature4Bias), .Out(data_11_array[j1][i1]));
    end
  endgenerate
  
  ////ROW 2
  generate
    localparam integer j2 = 2;
    for (i2 = 0; i2 < 24; i2 = i2 + 1)
    begin: addbit2
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j2+0][i2+0]), .Out(multi2[0][i2]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j2+0][i2+1]), .Out(multi2[1][i2]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j2+0][i2+2]), .Out(multi2[2][i2]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j2+0][i2+3]), .Out(multi2[3][i2]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j2+0][i2+4]), .Out(multi2[4][i2]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j2+1][i2+0]), .Out(multi2[5][i2]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j2+1][i2+1]), .Out(multi2[6][i2]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j2+1][i2+2]), .Out(multi2[7][i2]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j2+1][i2+3]), .Out(multi2[8][i2]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j2+1][i2+4]), .Out(multi2[9][i2]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j2+2][i2+0]), .Out(multi2[10][i2]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j2+2][i2+1]), .Out(multi2[11][i2]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j2+2][i2+2]), .Out(multi2[12][i2]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j2+2][i2+3]), .Out(multi2[13][i2]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j2+2][i2+4]), .Out(multi2[14][i2]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j2+3][i2+0]), .Out(multi2[15][i2]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j2+3][i2+1]), .Out(multi2[16][i2]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j2+3][i2+2]), .Out(multi2[17][i2]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j2+3][i2+3]), .Out(multi2[18][i2]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j2+3][i2+4]), .Out(multi2[19][i2]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j2+4][i2+0]), .Out(multi2[20][i2]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j2+4][i2+1]), .Out(multi2[21][i2]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j2+4][i2+2]), .Out(multi2[22][i2]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j2+4][i2+3]), .Out(multi2[23][i2]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j2+4][i2+4]), .Out(multi2[24][i2]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi2[0][i2]), .B(multi2[1][i2]), .Out(sum2[0][i2]));
      FP16_Add stage026(.A(multi2[2][i2]), .B(multi2[3][i2]), .Out(sum2[1][i2]));
      FP16_Add stage027(.A(multi2[4][i2]), .B(multi2[5][i2]), .Out(sum2[2][i2]));
      FP16_Add stage028(.A(multi2[6][i2]), .B(multi2[7][i2]), .Out(sum2[3][i2]));
      FP16_Add stage029(.A(multi2[8][i2]), .B(multi2[9][i2]), .Out(sum2[4][i2]));
      FP16_Add stage030(.A(multi2[10][i2]), .B(multi2[11][i2]), .Out(sum2[5][i2]));
      FP16_Add stage031(.A(multi2[12][i2]), .B(multi2[13][i2]), .Out(sum2[6][i2]));
      FP16_Add stage032(.A(multi2[14][i2]), .B(multi2[15][i2]), .Out(sum2[7][i2]));
      FP16_Add stage033(.A(multi2[16][i2]), .B(multi2[17][i2]), .Out(sum2[8][i2]));
      FP16_Add stage034(.A(multi2[18][i2]), .B(multi2[19][i2]), .Out(sum2[9][i2]));
      FP16_Add stage035(.A(multi2[20][i2]), .B(multi2[21][i2]), .Out(sum2[10][i2]));
      FP16_Add stage036(.A(multi2[22][i2]), .B(multi2[23][i2]), .Out(sum2[11][i2]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum2[0][i2]), .B(sum2[1][i2]), .Out(sum2[12][i2]));
      FP16_Add stage038(.A(sum2[2][i2]), .B(sum2[3][i2]), .Out(sum2[13][i2]));
      FP16_Add stage039(.A(sum2[4][i2]), .B(sum2[5][i2]), .Out(sum2[14][i2]));
      FP16_Add stage040(.A(sum2[6][i2]), .B(sum2[7][i2]), .Out(sum2[15][i2]));
      FP16_Add stage041(.A(sum2[8][i2]), .B(sum2[9][i2]), .Out(sum2[16][i2]));
      FP16_Add stage042(.A(sum2[10][i2]), .B(sum2[11][i2]), .Out(sum2[17][i2]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum2[12][i2]), .B(sum2[13][i2]), .Out(sum2[18][i2]));
      FP16_Add stage044(.A(sum2[14][i2]), .B(sum2[15][i2]), .Out(sum2[19][i2]));
      FP16_Add stage045(.A(sum2[16][i2]), .B(sum2[17][i2]), .Out(sum2[20][i2]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum2[18][i2]), .B(sum2[19][i2]), .Out(sum2[21][i2]));
      FP16_Add stage047(.A(sum2[20][i2]), .B(multi2[24][i2]), .Out(sum2[22][i2]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum2[21][i2]), .B(sum2[22][i2]), .Out(sum2[23][i2]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum2[23][i2]), .B(feature4Bias), .Out(data_11_array[j2][i2]));
    end
  endgenerate
  
  ////ROW 3
  generate
    localparam integer j3 = 3;
    for (i3 = 0; i3 < 24; i3 = i3 + 1)
    begin: addbit3
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j3+0][i3+0]), .Out(multi3[0][i3]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j3+0][i3+1]), .Out(multi3[1][i3]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j3+0][i3+2]), .Out(multi3[2][i3]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j3+0][i3+3]), .Out(multi3[3][i3]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j3+0][i3+4]), .Out(multi3[4][i3]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j3+1][i3+0]), .Out(multi3[5][i3]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j3+1][i3+1]), .Out(multi3[6][i3]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j3+1][i3+2]), .Out(multi3[7][i3]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j3+1][i3+3]), .Out(multi3[8][i3]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j3+1][i3+4]), .Out(multi3[9][i3]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j3+2][i3+0]), .Out(multi3[10][i3]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j3+2][i3+1]), .Out(multi3[11][i3]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j3+2][i3+2]), .Out(multi3[12][i3]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j3+2][i3+3]), .Out(multi3[13][i3]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j3+2][i3+4]), .Out(multi3[14][i3]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j3+3][i3+0]), .Out(multi3[15][i3]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j3+3][i3+1]), .Out(multi3[16][i3]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j3+3][i3+2]), .Out(multi3[17][i3]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j3+3][i3+3]), .Out(multi3[18][i3]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j3+3][i3+4]), .Out(multi3[19][i3]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j3+4][i3+0]), .Out(multi3[20][i3]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j3+4][i3+1]), .Out(multi3[21][i3]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j3+4][i3+2]), .Out(multi3[22][i3]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j3+4][i3+3]), .Out(multi3[23][i3]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j3+4][i3+4]), .Out(multi3[24][i3]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi3[0][i3]), .B(multi3[1][i3]), .Out(sum3[0][i3]));
      FP16_Add stage026(.A(multi3[2][i3]), .B(multi3[3][i3]), .Out(sum3[1][i3]));
      FP16_Add stage027(.A(multi3[4][i3]), .B(multi3[5][i3]), .Out(sum3[2][i3]));
      FP16_Add stage028(.A(multi3[6][i3]), .B(multi3[7][i3]), .Out(sum3[3][i3]));
      FP16_Add stage029(.A(multi3[8][i3]), .B(multi3[9][i3]), .Out(sum3[4][i3]));
      FP16_Add stage030(.A(multi3[10][i3]), .B(multi3[11][i3]), .Out(sum3[5][i3]));
      FP16_Add stage031(.A(multi3[12][i3]), .B(multi3[13][i3]), .Out(sum3[6][i3]));
      FP16_Add stage032(.A(multi3[14][i3]), .B(multi3[15][i3]), .Out(sum3[7][i3]));
      FP16_Add stage033(.A(multi3[16][i3]), .B(multi3[17][i3]), .Out(sum3[8][i3]));
      FP16_Add stage034(.A(multi3[18][i3]), .B(multi3[19][i3]), .Out(sum3[9][i3]));
      FP16_Add stage035(.A(multi3[20][i3]), .B(multi3[21][i3]), .Out(sum3[10][i3]));
      FP16_Add stage036(.A(multi3[22][i3]), .B(multi3[23][i3]), .Out(sum3[11][i3]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum3[0][i3]), .B(sum3[1][i3]), .Out(sum3[12][i3]));
      FP16_Add stage038(.A(sum3[2][i3]), .B(sum3[3][i3]), .Out(sum3[13][i3]));
      FP16_Add stage039(.A(sum3[4][i3]), .B(sum3[5][i3]), .Out(sum3[14][i3]));
      FP16_Add stage040(.A(sum3[6][i3]), .B(sum3[7][i3]), .Out(sum3[15][i3]));
      FP16_Add stage041(.A(sum3[8][i3]), .B(sum3[9][i3]), .Out(sum3[16][i3]));
      FP16_Add stage042(.A(sum3[10][i3]), .B(sum3[11][i3]), .Out(sum3[17][i3]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum3[12][i3]), .B(sum3[13][i3]), .Out(sum3[18][i3]));
      FP16_Add stage044(.A(sum3[14][i3]), .B(sum3[15][i3]), .Out(sum3[19][i3]));
      FP16_Add stage045(.A(sum3[16][i3]), .B(sum3[17][i3]), .Out(sum3[20][i3]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum3[18][i3]), .B(sum3[19][i3]), .Out(sum3[21][i3]));
      FP16_Add stage047(.A(sum3[20][i3]), .B(multi3[24][i3]), .Out(sum3[22][i3]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum3[21][i3]), .B(sum3[22][i3]), .Out(sum3[23][i3]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum3[23][i3]), .B(feature4Bias), .Out(data_11_array[j3][i3]));
    end
  endgenerate
  
  ////ROW 4
  generate
    localparam integer j4 = 4;
    for (i4 = 0; i4 < 24; i4 = i4 + 1)
    begin: addbit4
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j4+0][i4+0]), .Out(multi4[0][i4]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j4+0][i4+1]), .Out(multi4[1][i4]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j4+0][i4+2]), .Out(multi4[2][i4]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j4+0][i4+3]), .Out(multi4[3][i4]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j4+0][i4+4]), .Out(multi4[4][i4]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j4+1][i4+0]), .Out(multi4[5][i4]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j4+1][i4+1]), .Out(multi4[6][i4]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j4+1][i4+2]), .Out(multi4[7][i4]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j4+1][i4+3]), .Out(multi4[8][i4]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j4+1][i4+4]), .Out(multi4[9][i4]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j4+2][i4+0]), .Out(multi4[10][i4]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j4+2][i4+1]), .Out(multi4[11][i4]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j4+2][i4+2]), .Out(multi4[12][i4]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j4+2][i4+3]), .Out(multi4[13][i4]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j4+2][i4+4]), .Out(multi4[14][i4]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j4+3][i4+0]), .Out(multi4[15][i4]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j4+3][i4+1]), .Out(multi4[16][i4]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j4+3][i4+2]), .Out(multi4[17][i4]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j4+3][i4+3]), .Out(multi4[18][i4]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j4+3][i4+4]), .Out(multi4[19][i4]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j4+4][i4+0]), .Out(multi4[20][i4]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j4+4][i4+1]), .Out(multi4[21][i4]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j4+4][i4+2]), .Out(multi4[22][i4]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j4+4][i4+3]), .Out(multi4[23][i4]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j4+4][i4+4]), .Out(multi4[24][i4]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi4[0][i4]), .B(multi4[1][i4]), .Out(sum4[0][i4]));
      FP16_Add stage026(.A(multi4[2][i4]), .B(multi4[3][i4]), .Out(sum4[1][i4]));
      FP16_Add stage027(.A(multi4[4][i4]), .B(multi4[5][i4]), .Out(sum4[2][i4]));
      FP16_Add stage028(.A(multi4[6][i4]), .B(multi4[7][i4]), .Out(sum4[3][i4]));
      FP16_Add stage029(.A(multi4[8][i4]), .B(multi4[9][i4]), .Out(sum4[4][i4]));
      FP16_Add stage030(.A(multi4[10][i4]), .B(multi4[11][i4]), .Out(sum4[5][i4]));
      FP16_Add stage031(.A(multi4[12][i4]), .B(multi4[13][i4]), .Out(sum4[6][i4]));
      FP16_Add stage032(.A(multi4[14][i4]), .B(multi4[15][i4]), .Out(sum4[7][i4]));
      FP16_Add stage033(.A(multi4[16][i4]), .B(multi4[17][i4]), .Out(sum4[8][i4]));
      FP16_Add stage034(.A(multi4[18][i4]), .B(multi4[19][i4]), .Out(sum4[9][i4]));
      FP16_Add stage035(.A(multi4[20][i4]), .B(multi4[21][i4]), .Out(sum4[10][i4]));
      FP16_Add stage036(.A(multi4[22][i4]), .B(multi4[23][i4]), .Out(sum4[11][i4]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum4[0][i4]), .B(sum4[1][i4]), .Out(sum4[12][i4]));
      FP16_Add stage038(.A(sum4[2][i4]), .B(sum4[3][i4]), .Out(sum4[13][i4]));
      FP16_Add stage039(.A(sum4[4][i4]), .B(sum4[5][i4]), .Out(sum4[14][i4]));
      FP16_Add stage040(.A(sum4[6][i4]), .B(sum4[7][i4]), .Out(sum4[15][i4]));
      FP16_Add stage041(.A(sum4[8][i4]), .B(sum4[9][i4]), .Out(sum4[16][i4]));
      FP16_Add stage042(.A(sum4[10][i4]), .B(sum4[11][i4]), .Out(sum4[17][i4]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum4[12][i4]), .B(sum4[13][i4]), .Out(sum4[18][i4]));
      FP16_Add stage044(.A(sum4[14][i4]), .B(sum4[15][i4]), .Out(sum4[19][i4]));
      FP16_Add stage045(.A(sum4[16][i4]), .B(sum4[17][i4]), .Out(sum4[20][i4]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum4[18][i4]), .B(sum4[19][i4]), .Out(sum4[21][i4]));
      FP16_Add stage047(.A(sum4[20][i4]), .B(multi4[24][i4]), .Out(sum4[22][i4]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum4[21][i4]), .B(sum4[22][i4]), .Out(sum4[23][i4]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum4[23][i4]), .B(feature4Bias), .Out(data_11_array[j4][i4]));
    end
  endgenerate
  
  ////ROW 5
  generate
    localparam integer j5 = 5;
    for (i5 = 0; i5 < 24; i5 = i5 + 1)
    begin: addbit5
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j5+0][i5+0]), .Out(multi5[0][i5]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j5+0][i5+1]), .Out(multi5[1][i5]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j5+0][i5+2]), .Out(multi5[2][i5]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j5+0][i5+3]), .Out(multi5[3][i5]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j5+0][i5+4]), .Out(multi5[4][i5]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j5+1][i5+0]), .Out(multi5[5][i5]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j5+1][i5+1]), .Out(multi5[6][i5]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j5+1][i5+2]), .Out(multi5[7][i5]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j5+1][i5+3]), .Out(multi5[8][i5]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j5+1][i5+4]), .Out(multi5[9][i5]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j5+2][i5+0]), .Out(multi5[10][i5]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j5+2][i5+1]), .Out(multi5[11][i5]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j5+2][i5+2]), .Out(multi5[12][i5]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j5+2][i5+3]), .Out(multi5[13][i5]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j5+2][i5+4]), .Out(multi5[14][i5]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j5+3][i5+0]), .Out(multi5[15][i5]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j5+3][i5+1]), .Out(multi5[16][i5]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j5+3][i5+2]), .Out(multi5[17][i5]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j5+3][i5+3]), .Out(multi5[18][i5]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j5+3][i5+4]), .Out(multi5[19][i5]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j5+4][i5+0]), .Out(multi5[20][i5]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j5+4][i5+1]), .Out(multi5[21][i5]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j5+4][i5+2]), .Out(multi5[22][i5]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j5+4][i5+3]), .Out(multi5[23][i5]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j5+4][i5+4]), .Out(multi5[24][i5]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi5[0][i5]), .B(multi5[1][i5]), .Out(sum5[0][i5]));
      FP16_Add stage026(.A(multi5[2][i5]), .B(multi5[3][i5]), .Out(sum5[1][i5]));
      FP16_Add stage027(.A(multi5[4][i5]), .B(multi5[5][i5]), .Out(sum5[2][i5]));
      FP16_Add stage028(.A(multi5[6][i5]), .B(multi5[7][i5]), .Out(sum5[3][i5]));
      FP16_Add stage029(.A(multi5[8][i5]), .B(multi5[9][i5]), .Out(sum5[4][i5]));
      FP16_Add stage030(.A(multi5[10][i5]), .B(multi5[11][i5]), .Out(sum5[5][i5]));
      FP16_Add stage031(.A(multi5[12][i5]), .B(multi5[13][i5]), .Out(sum5[6][i5]));
      FP16_Add stage032(.A(multi5[14][i5]), .B(multi5[15][i5]), .Out(sum5[7][i5]));
      FP16_Add stage033(.A(multi5[16][i5]), .B(multi5[17][i5]), .Out(sum5[8][i5]));
      FP16_Add stage034(.A(multi5[18][i5]), .B(multi5[19][i5]), .Out(sum5[9][i5]));
      FP16_Add stage035(.A(multi5[20][i5]), .B(multi5[21][i5]), .Out(sum5[10][i5]));
      FP16_Add stage036(.A(multi5[22][i5]), .B(multi5[23][i5]), .Out(sum5[11][i5]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum5[0][i5]), .B(sum5[1][i5]), .Out(sum5[12][i5]));
      FP16_Add stage038(.A(sum5[2][i5]), .B(sum5[3][i5]), .Out(sum5[13][i5]));
      FP16_Add stage039(.A(sum5[4][i5]), .B(sum5[5][i5]), .Out(sum5[14][i5]));
      FP16_Add stage040(.A(sum5[6][i5]), .B(sum5[7][i5]), .Out(sum5[15][i5]));
      FP16_Add stage041(.A(sum5[8][i5]), .B(sum5[9][i5]), .Out(sum5[16][i5]));
      FP16_Add stage042(.A(sum5[10][i5]), .B(sum5[11][i5]), .Out(sum5[17][i5]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum5[12][i5]), .B(sum5[13][i5]), .Out(sum5[18][i5]));
      FP16_Add stage044(.A(sum5[14][i5]), .B(sum5[15][i5]), .Out(sum5[19][i5]));
      FP16_Add stage045(.A(sum5[16][i5]), .B(sum5[17][i5]), .Out(sum5[20][i5]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum5[18][i5]), .B(sum5[19][i5]), .Out(sum5[21][i5]));
      FP16_Add stage047(.A(sum5[20][i5]), .B(multi5[24][i5]), .Out(sum5[22][i5]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum5[21][i5]), .B(sum5[22][i5]), .Out(sum5[23][i5]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum5[23][i5]), .B(feature4Bias), .Out(data_11_array[j5][i5]));
    end
  endgenerate
  
  ////ROW 6
  generate
    localparam integer j6 = 6;
    for (i6 = 0; i6 < 24; i6 = i6 + 1)
    begin: addbit6
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j6+0][i6+0]), .Out(multi6[0][i6]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j6+0][i6+1]), .Out(multi6[1][i6]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j6+0][i6+2]), .Out(multi6[2][i6]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j6+0][i6+3]), .Out(multi6[3][i6]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j6+0][i6+4]), .Out(multi6[4][i6]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j6+1][i6+0]), .Out(multi6[5][i6]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j6+1][i6+1]), .Out(multi6[6][i6]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j6+1][i6+2]), .Out(multi6[7][i6]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j6+1][i6+3]), .Out(multi6[8][i6]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j6+1][i6+4]), .Out(multi6[9][i6]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j6+2][i6+0]), .Out(multi6[10][i6]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j6+2][i6+1]), .Out(multi6[11][i6]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j6+2][i6+2]), .Out(multi6[12][i6]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j6+2][i6+3]), .Out(multi6[13][i6]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j6+2][i6+4]), .Out(multi6[14][i6]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j6+3][i6+0]), .Out(multi6[15][i6]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j6+3][i6+1]), .Out(multi6[16][i6]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j6+3][i6+2]), .Out(multi6[17][i6]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j6+3][i6+3]), .Out(multi6[18][i6]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j6+3][i6+4]), .Out(multi6[19][i6]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j6+4][i6+0]), .Out(multi6[20][i6]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j6+4][i6+1]), .Out(multi6[21][i6]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j6+4][i6+2]), .Out(multi6[22][i6]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j6+4][i6+3]), .Out(multi6[23][i6]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j6+4][i6+4]), .Out(multi6[24][i6]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi6[0][i6]), .B(multi6[1][i6]), .Out(sum6[0][i6]));
      FP16_Add stage026(.A(multi6[2][i6]), .B(multi6[3][i6]), .Out(sum6[1][i6]));
      FP16_Add stage027(.A(multi6[4][i6]), .B(multi6[5][i6]), .Out(sum6[2][i6]));
      FP16_Add stage028(.A(multi6[6][i6]), .B(multi6[7][i6]), .Out(sum6[3][i6]));
      FP16_Add stage029(.A(multi6[8][i6]), .B(multi6[9][i6]), .Out(sum6[4][i6]));
      FP16_Add stage030(.A(multi6[10][i6]), .B(multi6[11][i6]), .Out(sum6[5][i6]));
      FP16_Add stage031(.A(multi6[12][i6]), .B(multi6[13][i6]), .Out(sum6[6][i6]));
      FP16_Add stage032(.A(multi6[14][i6]), .B(multi6[15][i6]), .Out(sum6[7][i6]));
      FP16_Add stage033(.A(multi6[16][i6]), .B(multi6[17][i6]), .Out(sum6[8][i6]));
      FP16_Add stage034(.A(multi6[18][i6]), .B(multi6[19][i6]), .Out(sum6[9][i6]));
      FP16_Add stage035(.A(multi6[20][i6]), .B(multi6[21][i6]), .Out(sum6[10][i6]));
      FP16_Add stage036(.A(multi6[22][i6]), .B(multi6[23][i6]), .Out(sum6[11][i6]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum6[0][i6]), .B(sum6[1][i6]), .Out(sum6[12][i6]));
      FP16_Add stage038(.A(sum6[2][i6]), .B(sum6[3][i6]), .Out(sum6[13][i6]));
      FP16_Add stage039(.A(sum6[4][i6]), .B(sum6[5][i6]), .Out(sum6[14][i6]));
      FP16_Add stage040(.A(sum6[6][i6]), .B(sum6[7][i6]), .Out(sum6[15][i6]));
      FP16_Add stage041(.A(sum6[8][i6]), .B(sum6[9][i6]), .Out(sum6[16][i6]));
      FP16_Add stage042(.A(sum6[10][i6]), .B(sum6[11][i6]), .Out(sum6[17][i6]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum6[12][i6]), .B(sum6[13][i6]), .Out(sum6[18][i6]));
      FP16_Add stage044(.A(sum6[14][i6]), .B(sum6[15][i6]), .Out(sum6[19][i6]));
      FP16_Add stage045(.A(sum6[16][i6]), .B(sum6[17][i6]), .Out(sum6[20][i6]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum6[18][i6]), .B(sum6[19][i6]), .Out(sum6[21][i6]));
      FP16_Add stage047(.A(sum6[20][i6]), .B(multi6[24][i6]), .Out(sum6[22][i6]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum6[21][i6]), .B(sum6[22][i6]), .Out(sum6[23][i6]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum6[23][i6]), .B(feature4Bias), .Out(data_11_array[j6][i6]));
    end
  endgenerate
  
  ////ROW 7
  generate
    localparam integer j7 = 7;
    for (i7 = 0; i7 < 24; i7 = i7 + 1)
    begin: addbit7
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j7+0][i7+0]), .Out(multi7[0][i7]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j7+0][i7+1]), .Out(multi7[1][i7]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j7+0][i7+2]), .Out(multi7[2][i7]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j7+0][i7+3]), .Out(multi7[3][i7]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j7+0][i7+4]), .Out(multi7[4][i7]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j7+1][i7+0]), .Out(multi7[5][i7]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j7+1][i7+1]), .Out(multi7[6][i7]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j7+1][i7+2]), .Out(multi7[7][i7]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j7+1][i7+3]), .Out(multi7[8][i7]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j7+1][i7+4]), .Out(multi7[9][i7]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j7+2][i7+0]), .Out(multi7[10][i7]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j7+2][i7+1]), .Out(multi7[11][i7]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j7+2][i7+2]), .Out(multi7[12][i7]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j7+2][i7+3]), .Out(multi7[13][i7]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j7+2][i7+4]), .Out(multi7[14][i7]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j7+3][i7+0]), .Out(multi7[15][i7]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j7+3][i7+1]), .Out(multi7[16][i7]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j7+3][i7+2]), .Out(multi7[17][i7]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j7+3][i7+3]), .Out(multi7[18][i7]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j7+3][i7+4]), .Out(multi7[19][i7]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j7+4][i7+0]), .Out(multi7[20][i7]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j7+4][i7+1]), .Out(multi7[21][i7]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j7+4][i7+2]), .Out(multi7[22][i7]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j7+4][i7+3]), .Out(multi7[23][i7]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j7+4][i7+4]), .Out(multi7[24][i7]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi7[0][i7]), .B(multi7[1][i7]), .Out(sum7[0][i7]));
      FP16_Add stage026(.A(multi7[2][i7]), .B(multi7[3][i7]), .Out(sum7[1][i7]));
      FP16_Add stage027(.A(multi7[4][i7]), .B(multi7[5][i7]), .Out(sum7[2][i7]));
      FP16_Add stage028(.A(multi7[6][i7]), .B(multi7[7][i7]), .Out(sum7[3][i7]));
      FP16_Add stage029(.A(multi7[8][i7]), .B(multi7[9][i7]), .Out(sum7[4][i7]));
      FP16_Add stage030(.A(multi7[10][i7]), .B(multi7[11][i7]), .Out(sum7[5][i7]));
      FP16_Add stage031(.A(multi7[12][i7]), .B(multi7[13][i7]), .Out(sum7[6][i7]));
      FP16_Add stage032(.A(multi7[14][i7]), .B(multi7[15][i7]), .Out(sum7[7][i7]));
      FP16_Add stage033(.A(multi7[16][i7]), .B(multi7[17][i7]), .Out(sum7[8][i7]));
      FP16_Add stage034(.A(multi7[18][i7]), .B(multi7[19][i7]), .Out(sum7[9][i7]));
      FP16_Add stage035(.A(multi7[20][i7]), .B(multi7[21][i7]), .Out(sum7[10][i7]));
      FP16_Add stage036(.A(multi7[22][i7]), .B(multi7[23][i7]), .Out(sum7[11][i7]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum7[0][i7]), .B(sum7[1][i7]), .Out(sum7[12][i7]));
      FP16_Add stage038(.A(sum7[2][i7]), .B(sum7[3][i7]), .Out(sum7[13][i7]));
      FP16_Add stage039(.A(sum7[4][i7]), .B(sum7[5][i7]), .Out(sum7[14][i7]));
      FP16_Add stage040(.A(sum7[6][i7]), .B(sum7[7][i7]), .Out(sum7[15][i7]));
      FP16_Add stage041(.A(sum7[8][i7]), .B(sum7[9][i7]), .Out(sum7[16][i7]));
      FP16_Add stage042(.A(sum7[10][i7]), .B(sum7[11][i7]), .Out(sum7[17][i7]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum7[12][i7]), .B(sum7[13][i7]), .Out(sum7[18][i7]));
      FP16_Add stage044(.A(sum7[14][i7]), .B(sum7[15][i7]), .Out(sum7[19][i7]));
      FP16_Add stage045(.A(sum7[16][i7]), .B(sum7[17][i7]), .Out(sum7[20][i7]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum7[18][i7]), .B(sum7[19][i7]), .Out(sum7[21][i7]));
      FP16_Add stage047(.A(sum7[20][i7]), .B(multi7[24][i7]), .Out(sum7[22][i7]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum7[21][i7]), .B(sum7[22][i7]), .Out(sum7[23][i7]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum7[23][i7]), .B(feature4Bias), .Out(data_11_array[j7][i7]));
    end
  endgenerate
  
  ////ROW 8
  generate
    localparam integer j8 = 8;
    for (i8 = 0; i8 < 24; i8 = i8 + 1)
    begin: addbit8
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j8+0][i8+0]), .Out(multi8[0][i8]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j8+0][i8+1]), .Out(multi8[1][i8]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j8+0][i8+2]), .Out(multi8[2][i8]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j8+0][i8+3]), .Out(multi8[3][i8]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j8+0][i8+4]), .Out(multi8[4][i8]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j8+1][i8+0]), .Out(multi8[5][i8]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j8+1][i8+1]), .Out(multi8[6][i8]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j8+1][i8+2]), .Out(multi8[7][i8]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j8+1][i8+3]), .Out(multi8[8][i8]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j8+1][i8+4]), .Out(multi8[9][i8]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j8+2][i8+0]), .Out(multi8[10][i8]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j8+2][i8+1]), .Out(multi8[11][i8]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j8+2][i8+2]), .Out(multi8[12][i8]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j8+2][i8+3]), .Out(multi8[13][i8]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j8+2][i8+4]), .Out(multi8[14][i8]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j8+3][i8+0]), .Out(multi8[15][i8]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j8+3][i8+1]), .Out(multi8[16][i8]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j8+3][i8+2]), .Out(multi8[17][i8]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j8+3][i8+3]), .Out(multi8[18][i8]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j8+3][i8+4]), .Out(multi8[19][i8]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j8+4][i8+0]), .Out(multi8[20][i8]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j8+4][i8+1]), .Out(multi8[21][i8]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j8+4][i8+2]), .Out(multi8[22][i8]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j8+4][i8+3]), .Out(multi8[23][i8]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j8+4][i8+4]), .Out(multi8[24][i8]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi8[0][i8]), .B(multi8[1][i8]), .Out(sum8[0][i8]));
      FP16_Add stage026(.A(multi8[2][i8]), .B(multi8[3][i8]), .Out(sum8[1][i8]));
      FP16_Add stage027(.A(multi8[4][i8]), .B(multi8[5][i8]), .Out(sum8[2][i8]));
      FP16_Add stage028(.A(multi8[6][i8]), .B(multi8[7][i8]), .Out(sum8[3][i8]));
      FP16_Add stage029(.A(multi8[8][i8]), .B(multi8[9][i8]), .Out(sum8[4][i8]));
      FP16_Add stage030(.A(multi8[10][i8]), .B(multi8[11][i8]), .Out(sum8[5][i8]));
      FP16_Add stage031(.A(multi8[12][i8]), .B(multi8[13][i8]), .Out(sum8[6][i8]));
      FP16_Add stage032(.A(multi8[14][i8]), .B(multi8[15][i8]), .Out(sum8[7][i8]));
      FP16_Add stage033(.A(multi8[16][i8]), .B(multi8[17][i8]), .Out(sum8[8][i8]));
      FP16_Add stage034(.A(multi8[18][i8]), .B(multi8[19][i8]), .Out(sum8[9][i8]));
      FP16_Add stage035(.A(multi8[20][i8]), .B(multi8[21][i8]), .Out(sum8[10][i8]));
      FP16_Add stage036(.A(multi8[22][i8]), .B(multi8[23][i8]), .Out(sum8[11][i8]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum8[0][i8]), .B(sum8[1][i8]), .Out(sum8[12][i8]));
      FP16_Add stage038(.A(sum8[2][i8]), .B(sum8[3][i8]), .Out(sum8[13][i8]));
      FP16_Add stage039(.A(sum8[4][i8]), .B(sum8[5][i8]), .Out(sum8[14][i8]));
      FP16_Add stage040(.A(sum8[6][i8]), .B(sum8[7][i8]), .Out(sum8[15][i8]));
      FP16_Add stage041(.A(sum8[8][i8]), .B(sum8[9][i8]), .Out(sum8[16][i8]));
      FP16_Add stage042(.A(sum8[10][i8]), .B(sum8[11][i8]), .Out(sum8[17][i8]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum8[12][i8]), .B(sum8[13][i8]), .Out(sum8[18][i8]));
      FP16_Add stage044(.A(sum8[14][i8]), .B(sum8[15][i8]), .Out(sum8[19][i8]));
      FP16_Add stage045(.A(sum8[16][i8]), .B(sum8[17][i8]), .Out(sum8[20][i8]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum8[18][i8]), .B(sum8[19][i8]), .Out(sum8[21][i8]));
      FP16_Add stage047(.A(sum8[20][i8]), .B(multi8[24][i8]), .Out(sum8[22][i8]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum8[21][i8]), .B(sum8[22][i8]), .Out(sum8[23][i8]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum8[23][i8]), .B(feature4Bias), .Out(data_11_array[j8][i8]));
    end
  endgenerate
  
  ////ROW 9
  generate
    localparam integer j9 = 9;
    for (i9 = 0; i9 < 24; i9 = i9 + 1)
    begin: addbit9
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j9+0][i9+0]), .Out(multi9[0][i9]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j9+0][i9+1]), .Out(multi9[1][i9]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j9+0][i9+2]), .Out(multi9[2][i9]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j9+0][i9+3]), .Out(multi9[3][i9]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j9+0][i9+4]), .Out(multi9[4][i9]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j9+1][i9+0]), .Out(multi9[5][i9]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j9+1][i9+1]), .Out(multi9[6][i9]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j9+1][i9+2]), .Out(multi9[7][i9]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j9+1][i9+3]), .Out(multi9[8][i9]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j9+1][i9+4]), .Out(multi9[9][i9]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j9+2][i9+0]), .Out(multi9[10][i9]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j9+2][i9+1]), .Out(multi9[11][i9]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j9+2][i9+2]), .Out(multi9[12][i9]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j9+2][i9+3]), .Out(multi9[13][i9]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j9+2][i9+4]), .Out(multi9[14][i9]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j9+3][i9+0]), .Out(multi9[15][i9]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j9+3][i9+1]), .Out(multi9[16][i9]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j9+3][i9+2]), .Out(multi9[17][i9]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j9+3][i9+3]), .Out(multi9[18][i9]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j9+3][i9+4]), .Out(multi9[19][i9]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j9+4][i9+0]), .Out(multi9[20][i9]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j9+4][i9+1]), .Out(multi9[21][i9]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j9+4][i9+2]), .Out(multi9[22][i9]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j9+4][i9+3]), .Out(multi9[23][i9]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j9+4][i9+4]), .Out(multi9[24][i9]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi9[0][i9]), .B(multi9[1][i9]), .Out(sum9[0][i9]));
      FP16_Add stage026(.A(multi9[2][i9]), .B(multi9[3][i9]), .Out(sum9[1][i9]));
      FP16_Add stage027(.A(multi9[4][i9]), .B(multi9[5][i9]), .Out(sum9[2][i9]));
      FP16_Add stage028(.A(multi9[6][i9]), .B(multi9[7][i9]), .Out(sum9[3][i9]));
      FP16_Add stage029(.A(multi9[8][i9]), .B(multi9[9][i9]), .Out(sum9[4][i9]));
      FP16_Add stage030(.A(multi9[10][i9]), .B(multi9[11][i9]), .Out(sum9[5][i9]));
      FP16_Add stage031(.A(multi9[12][i9]), .B(multi9[13][i9]), .Out(sum9[6][i9]));
      FP16_Add stage032(.A(multi9[14][i9]), .B(multi9[15][i9]), .Out(sum9[7][i9]));
      FP16_Add stage033(.A(multi9[16][i9]), .B(multi9[17][i9]), .Out(sum9[8][i9]));
      FP16_Add stage034(.A(multi9[18][i9]), .B(multi9[19][i9]), .Out(sum9[9][i9]));
      FP16_Add stage035(.A(multi9[20][i9]), .B(multi9[21][i9]), .Out(sum9[10][i9]));
      FP16_Add stage036(.A(multi9[22][i9]), .B(multi9[23][i9]), .Out(sum9[11][i9]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum9[0][i9]), .B(sum9[1][i9]), .Out(sum9[12][i9]));
      FP16_Add stage038(.A(sum9[2][i9]), .B(sum9[3][i9]), .Out(sum9[13][i9]));
      FP16_Add stage039(.A(sum9[4][i9]), .B(sum9[5][i9]), .Out(sum9[14][i9]));
      FP16_Add stage040(.A(sum9[6][i9]), .B(sum9[7][i9]), .Out(sum9[15][i9]));
      FP16_Add stage041(.A(sum9[8][i9]), .B(sum9[9][i9]), .Out(sum9[16][i9]));
      FP16_Add stage042(.A(sum9[10][i9]), .B(sum9[11][i9]), .Out(sum9[17][i9]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum9[12][i9]), .B(sum9[13][i9]), .Out(sum9[18][i9]));
      FP16_Add stage044(.A(sum9[14][i9]), .B(sum9[15][i9]), .Out(sum9[19][i9]));
      FP16_Add stage045(.A(sum9[16][i9]), .B(sum9[17][i9]), .Out(sum9[20][i9]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum9[18][i9]), .B(sum9[19][i9]), .Out(sum9[21][i9]));
      FP16_Add stage047(.A(sum9[20][i9]), .B(multi9[24][i9]), .Out(sum9[22][i9]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum9[21][i9]), .B(sum9[22][i9]), .Out(sum9[23][i9]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum9[23][i9]), .B(feature4Bias), .Out(data_11_array[j9][i9]));
    end
  endgenerate
  
  ////ROW 10
  generate
    localparam integer j10 = 10;
    for (i10 = 0; i10 < 24; i10 = i10 + 1)
    begin: addbit10
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j10+0][i10+0]), .Out(multi10[0][i10]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j10+0][i10+1]), .Out(multi10[1][i10]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j10+0][i10+2]), .Out(multi10[2][i10]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j10+0][i10+3]), .Out(multi10[3][i10]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j10+0][i10+4]), .Out(multi10[4][i10]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j10+1][i10+0]), .Out(multi10[5][i10]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j10+1][i10+1]), .Out(multi10[6][i10]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j10+1][i10+2]), .Out(multi10[7][i10]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j10+1][i10+3]), .Out(multi10[8][i10]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j10+1][i10+4]), .Out(multi10[9][i10]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j10+2][i10+0]), .Out(multi10[10][i10]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j10+2][i10+1]), .Out(multi10[11][i10]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j10+2][i10+2]), .Out(multi10[12][i10]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j10+2][i10+3]), .Out(multi10[13][i10]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j10+2][i10+4]), .Out(multi10[14][i10]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j10+3][i10+0]), .Out(multi10[15][i10]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j10+3][i10+1]), .Out(multi10[16][i10]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j10+3][i10+2]), .Out(multi10[17][i10]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j10+3][i10+3]), .Out(multi10[18][i10]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j10+3][i10+4]), .Out(multi10[19][i10]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j10+4][i10+0]), .Out(multi10[20][i10]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j10+4][i10+1]), .Out(multi10[21][i10]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j10+4][i10+2]), .Out(multi10[22][i10]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j10+4][i10+3]), .Out(multi10[23][i10]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j10+4][i10+4]), .Out(multi10[24][i10]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi10[0][i10]), .B(multi10[1][i10]), .Out(sum10[0][i10]));
      FP16_Add stage026(.A(multi10[2][i10]), .B(multi10[3][i10]), .Out(sum10[1][i10]));
      FP16_Add stage027(.A(multi10[4][i10]), .B(multi10[5][i10]), .Out(sum10[2][i10]));
      FP16_Add stage028(.A(multi10[6][i10]), .B(multi10[7][i10]), .Out(sum10[3][i10]));
      FP16_Add stage029(.A(multi10[8][i10]), .B(multi10[9][i10]), .Out(sum10[4][i10]));
      FP16_Add stage030(.A(multi10[10][i10]), .B(multi10[11][i10]), .Out(sum10[5][i10]));
      FP16_Add stage031(.A(multi10[12][i10]), .B(multi10[13][i10]), .Out(sum10[6][i10]));
      FP16_Add stage032(.A(multi10[14][i10]), .B(multi10[15][i10]), .Out(sum10[7][i10]));
      FP16_Add stage033(.A(multi10[16][i10]), .B(multi10[17][i10]), .Out(sum10[8][i10]));
      FP16_Add stage034(.A(multi10[18][i10]), .B(multi10[19][i10]), .Out(sum10[9][i10]));
      FP16_Add stage035(.A(multi10[20][i10]), .B(multi10[21][i10]), .Out(sum10[10][i10]));
      FP16_Add stage036(.A(multi10[22][i10]), .B(multi10[23][i10]), .Out(sum10[11][i10]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum10[0][i10]), .B(sum10[1][i10]), .Out(sum10[12][i10]));
      FP16_Add stage038(.A(sum10[2][i10]), .B(sum10[3][i10]), .Out(sum10[13][i10]));
      FP16_Add stage039(.A(sum10[4][i10]), .B(sum10[5][i10]), .Out(sum10[14][i10]));
      FP16_Add stage040(.A(sum10[6][i10]), .B(sum10[7][i10]), .Out(sum10[15][i10]));
      FP16_Add stage041(.A(sum10[8][i10]), .B(sum10[9][i10]), .Out(sum10[16][i10]));
      FP16_Add stage042(.A(sum10[10][i10]), .B(sum10[11][i10]), .Out(sum10[17][i10]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum10[12][i10]), .B(sum10[13][i10]), .Out(sum10[18][i10]));
      FP16_Add stage044(.A(sum10[14][i10]), .B(sum10[15][i10]), .Out(sum10[19][i10]));
      FP16_Add stage045(.A(sum10[16][i10]), .B(sum10[17][i10]), .Out(sum10[20][i10]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum10[18][i10]), .B(sum10[19][i10]), .Out(sum10[21][i10]));
      FP16_Add stage047(.A(sum10[20][i10]), .B(multi10[24][i10]), .Out(sum10[22][i10]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum10[21][i10]), .B(sum10[22][i10]), .Out(sum10[23][i10]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum10[23][i10]), .B(feature4Bias), .Out(data_11_array[j10][i10]));
    end
  endgenerate
  
    ////ROW 11
  generate
    localparam integer j11 = 11;
    for (i11 = 0; i11 < 24; i11 = i11 + 1)
    begin: addbit11
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j11+0][i11+0]), .Out(multi11[0][i11]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j11+0][i11+1]), .Out(multi11[1][i11]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j11+0][i11+2]), .Out(multi11[2][i11]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j11+0][i11+3]), .Out(multi11[3][i11]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j11+0][i11+4]), .Out(multi11[4][i11]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j11+1][i11+0]), .Out(multi11[5][i11]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j11+1][i11+1]), .Out(multi11[6][i11]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j11+1][i11+2]), .Out(multi11[7][i11]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j11+1][i11+3]), .Out(multi11[8][i11]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j11+1][i11+4]), .Out(multi11[9][i11]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j11+2][i11+0]), .Out(multi11[10][i11]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j11+2][i11+1]), .Out(multi11[11][i11]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j11+2][i11+2]), .Out(multi11[12][i11]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j11+2][i11+3]), .Out(multi11[13][i11]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j11+2][i11+4]), .Out(multi11[14][i11]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j11+3][i11+0]), .Out(multi11[15][i11]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j11+3][i11+1]), .Out(multi11[16][i11]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j11+3][i11+2]), .Out(multi11[17][i11]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j11+3][i11+3]), .Out(multi11[18][i11]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j11+3][i11+4]), .Out(multi11[19][i11]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j11+4][i11+0]), .Out(multi11[20][i11]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j11+4][i11+1]), .Out(multi11[21][i11]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j11+4][i11+2]), .Out(multi11[22][i11]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j11+4][i11+3]), .Out(multi11[23][i11]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j11+4][i11+4]), .Out(multi11[24][i11]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi11[0][i11]), .B(multi11[1][i11]), .Out(sum11[0][i11]));
      FP16_Add stage026(.A(multi11[2][i11]), .B(multi11[3][i11]), .Out(sum11[1][i11]));
      FP16_Add stage027(.A(multi11[4][i11]), .B(multi11[5][i11]), .Out(sum11[2][i11]));
      FP16_Add stage028(.A(multi11[6][i11]), .B(multi11[7][i11]), .Out(sum11[3][i11]));
      FP16_Add stage029(.A(multi11[8][i11]), .B(multi11[9][i11]), .Out(sum11[4][i11]));
      FP16_Add stage030(.A(multi11[10][i11]), .B(multi11[11][i11]), .Out(sum11[5][i11]));
      FP16_Add stage031(.A(multi11[12][i11]), .B(multi11[13][i11]), .Out(sum11[6][i11]));
      FP16_Add stage032(.A(multi11[14][i11]), .B(multi11[15][i11]), .Out(sum11[7][i11]));
      FP16_Add stage033(.A(multi11[16][i11]), .B(multi11[17][i11]), .Out(sum11[8][i11]));
      FP16_Add stage034(.A(multi11[18][i11]), .B(multi11[19][i11]), .Out(sum11[9][i11]));
      FP16_Add stage035(.A(multi11[20][i11]), .B(multi11[21][i11]), .Out(sum11[10][i11]));
      FP16_Add stage036(.A(multi11[22][i11]), .B(multi11[23][i11]), .Out(sum11[11][i11]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum11[0][i11]), .B(sum11[1][i11]), .Out(sum11[12][i11]));
      FP16_Add stage038(.A(sum11[2][i11]), .B(sum11[3][i11]), .Out(sum11[13][i11]));
      FP16_Add stage039(.A(sum11[4][i11]), .B(sum11[5][i11]), .Out(sum11[14][i11]));
      FP16_Add stage040(.A(sum11[6][i11]), .B(sum11[7][i11]), .Out(sum11[15][i11]));
      FP16_Add stage041(.A(sum11[8][i11]), .B(sum11[9][i11]), .Out(sum11[16][i11]));
      FP16_Add stage042(.A(sum11[10][i11]), .B(sum11[11][i11]), .Out(sum11[17][i11]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum11[12][i11]), .B(sum11[13][i11]), .Out(sum11[18][i11]));
      FP16_Add stage044(.A(sum11[14][i11]), .B(sum11[15][i11]), .Out(sum11[19][i11]));
      FP16_Add stage045(.A(sum11[16][i11]), .B(sum11[17][i11]), .Out(sum11[20][i11]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum11[18][i11]), .B(sum11[19][i11]), .Out(sum11[21][i11]));
      FP16_Add stage047(.A(sum11[20][i11]), .B(multi11[24][i11]), .Out(sum11[22][i11]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum11[21][i11]), .B(sum11[22][i11]), .Out(sum11[23][i11]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum11[23][i11]), .B(feature4Bias), .Out(data_11_array[j11][i11]));
    end
  endgenerate

  ////ROW 12
  generate
    localparam integer j12 = 12;
    for (i12 = 0; i12 < 24; i12 = i12 + 1)
    begin: addbit12
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j12+0][i12+0]), .Out(multi12[0][i12]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j12+0][i12+1]), .Out(multi12[1][i12]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j12+0][i12+2]), .Out(multi12[2][i12]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j12+0][i12+3]), .Out(multi12[3][i12]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j12+0][i12+4]), .Out(multi12[4][i12]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j12+1][i12+0]), .Out(multi12[5][i12]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j12+1][i12+1]), .Out(multi12[6][i12]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j12+1][i12+2]), .Out(multi12[7][i12]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j12+1][i12+3]), .Out(multi12[8][i12]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j12+1][i12+4]), .Out(multi12[9][i12]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j12+2][i12+0]), .Out(multi12[10][i12]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j12+2][i12+1]), .Out(multi12[11][i12]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j12+2][i12+2]), .Out(multi12[12][i12]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j12+2][i12+3]), .Out(multi12[13][i12]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j12+2][i12+4]), .Out(multi12[14][i12]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j12+3][i12+0]), .Out(multi12[15][i12]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j12+3][i12+1]), .Out(multi12[16][i12]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j12+3][i12+2]), .Out(multi12[17][i12]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j12+3][i12+3]), .Out(multi12[18][i12]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j12+3][i12+4]), .Out(multi12[19][i12]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j12+4][i12+0]), .Out(multi12[20][i12]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j12+4][i12+1]), .Out(multi12[21][i12]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j12+4][i12+2]), .Out(multi12[22][i12]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j12+4][i12+3]), .Out(multi12[23][i12]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j12+4][i12+4]), .Out(multi12[24][i12]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi12[0][i12]), .B(multi12[1][i12]), .Out(sum12[0][i12]));
      FP16_Add stage026(.A(multi12[2][i12]), .B(multi12[3][i12]), .Out(sum12[1][i12]));
      FP16_Add stage027(.A(multi12[4][i12]), .B(multi12[5][i12]), .Out(sum12[2][i12]));
      FP16_Add stage028(.A(multi12[6][i12]), .B(multi12[7][i12]), .Out(sum12[3][i12]));
      FP16_Add stage029(.A(multi12[8][i12]), .B(multi12[9][i12]), .Out(sum12[4][i12]));
      FP16_Add stage030(.A(multi12[10][i12]), .B(multi12[11][i12]), .Out(sum12[5][i12]));
      FP16_Add stage031(.A(multi12[12][i12]), .B(multi12[13][i12]), .Out(sum12[6][i12]));
      FP16_Add stage032(.A(multi12[14][i12]), .B(multi12[15][i12]), .Out(sum12[7][i12]));
      FP16_Add stage033(.A(multi12[16][i12]), .B(multi12[17][i12]), .Out(sum12[8][i12]));
      FP16_Add stage034(.A(multi12[18][i12]), .B(multi12[19][i12]), .Out(sum12[9][i12]));
      FP16_Add stage035(.A(multi12[20][i12]), .B(multi12[21][i12]), .Out(sum12[10][i12]));
      FP16_Add stage036(.A(multi12[22][i12]), .B(multi12[23][i12]), .Out(sum12[11][i12]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum12[0][i12]), .B(sum12[1][i12]), .Out(sum12[12][i12]));
      FP16_Add stage038(.A(sum12[2][i12]), .B(sum12[3][i12]), .Out(sum12[13][i12]));
      FP16_Add stage039(.A(sum12[4][i12]), .B(sum12[5][i12]), .Out(sum12[14][i12]));
      FP16_Add stage040(.A(sum12[6][i12]), .B(sum12[7][i12]), .Out(sum12[15][i12]));
      FP16_Add stage041(.A(sum12[8][i12]), .B(sum12[9][i12]), .Out(sum12[16][i12]));
      FP16_Add stage042(.A(sum12[10][i12]), .B(sum12[11][i12]), .Out(sum12[17][i12]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum12[12][i12]), .B(sum12[13][i12]), .Out(sum12[18][i12]));
      FP16_Add stage044(.A(sum12[14][i12]), .B(sum12[15][i12]), .Out(sum12[19][i12]));
      FP16_Add stage045(.A(sum12[16][i12]), .B(sum12[17][i12]), .Out(sum12[20][i12]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum12[18][i12]), .B(sum12[19][i12]), .Out(sum12[21][i12]));
      FP16_Add stage047(.A(sum12[20][i12]), .B(multi12[24][i12]), .Out(sum12[22][i12]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum12[21][i12]), .B(sum12[22][i12]), .Out(sum12[23][i12]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum12[23][i12]), .B(feature4Bias), .Out(data_11_array[j12][i12]));
    end
  endgenerate

  ////ROW 13
  generate
    localparam integer j13 = 13;
    for (i13 = 0; i13 < 24; i13 = i13 + 1)
    begin: addbit13
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j13+0][i13+0]), .Out(multi13[0][i13]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j13+0][i13+1]), .Out(multi13[1][i13]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j13+0][i13+2]), .Out(multi13[2][i13]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j13+0][i13+3]), .Out(multi13[3][i13]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j13+0][i13+4]), .Out(multi13[4][i13]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j13+1][i13+0]), .Out(multi13[5][i13]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j13+1][i13+1]), .Out(multi13[6][i13]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j13+1][i13+2]), .Out(multi13[7][i13]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j13+1][i13+3]), .Out(multi13[8][i13]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j13+1][i13+4]), .Out(multi13[9][i13]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j13+2][i13+0]), .Out(multi13[10][i13]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j13+2][i13+1]), .Out(multi13[11][i13]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j13+2][i13+2]), .Out(multi13[12][i13]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j13+2][i13+3]), .Out(multi13[13][i13]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j13+2][i13+4]), .Out(multi13[14][i13]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j13+3][i13+0]), .Out(multi13[15][i13]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j13+3][i13+1]), .Out(multi13[16][i13]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j13+3][i13+2]), .Out(multi13[17][i13]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j13+3][i13+3]), .Out(multi13[18][i13]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j13+3][i13+4]), .Out(multi13[19][i13]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j13+4][i13+0]), .Out(multi13[20][i13]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j13+4][i13+1]), .Out(multi13[21][i13]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j13+4][i13+2]), .Out(multi13[22][i13]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j13+4][i13+3]), .Out(multi13[23][i13]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j13+4][i13+4]), .Out(multi13[24][i13]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi13[0][i13]), .B(multi13[1][i13]), .Out(sum13[0][i13]));
      FP16_Add stage026(.A(multi13[2][i13]), .B(multi13[3][i13]), .Out(sum13[1][i13]));
      FP16_Add stage027(.A(multi13[4][i13]), .B(multi13[5][i13]), .Out(sum13[2][i13]));
      FP16_Add stage028(.A(multi13[6][i13]), .B(multi13[7][i13]), .Out(sum13[3][i13]));
      FP16_Add stage029(.A(multi13[8][i13]), .B(multi13[9][i13]), .Out(sum13[4][i13]));
      FP16_Add stage030(.A(multi13[10][i13]), .B(multi13[11][i13]), .Out(sum13[5][i13]));
      FP16_Add stage031(.A(multi13[12][i13]), .B(multi13[13][i13]), .Out(sum13[6][i13]));
      FP16_Add stage032(.A(multi13[14][i13]), .B(multi13[15][i13]), .Out(sum13[7][i13]));
      FP16_Add stage033(.A(multi13[16][i13]), .B(multi13[17][i13]), .Out(sum13[8][i13]));
      FP16_Add stage034(.A(multi13[18][i13]), .B(multi13[19][i13]), .Out(sum13[9][i13]));
      FP16_Add stage035(.A(multi13[20][i13]), .B(multi13[21][i13]), .Out(sum13[10][i13]));
      FP16_Add stage036(.A(multi13[22][i13]), .B(multi13[23][i13]), .Out(sum13[11][i13]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum13[0][i13]), .B(sum13[1][i13]), .Out(sum13[12][i13]));
      FP16_Add stage038(.A(sum13[2][i13]), .B(sum13[3][i13]), .Out(sum13[13][i13]));
      FP16_Add stage039(.A(sum13[4][i13]), .B(sum13[5][i13]), .Out(sum13[14][i13]));
      FP16_Add stage040(.A(sum13[6][i13]), .B(sum13[7][i13]), .Out(sum13[15][i13]));
      FP16_Add stage041(.A(sum13[8][i13]), .B(sum13[9][i13]), .Out(sum13[16][i13]));
      FP16_Add stage042(.A(sum13[10][i13]), .B(sum13[11][i13]), .Out(sum13[17][i13]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum13[12][i13]), .B(sum13[13][i13]), .Out(sum13[18][i13]));
      FP16_Add stage044(.A(sum13[14][i13]), .B(sum13[15][i13]), .Out(sum13[19][i13]));
      FP16_Add stage045(.A(sum13[16][i13]), .B(sum13[17][i13]), .Out(sum13[20][i13]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum13[18][i13]), .B(sum13[19][i13]), .Out(sum13[21][i13]));
      FP16_Add stage047(.A(sum13[20][i13]), .B(multi13[24][i13]), .Out(sum13[22][i13]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum13[21][i13]), .B(sum13[22][i13]), .Out(sum13[23][i13]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum13[23][i13]), .B(feature4Bias), .Out(data_11_array[j13][i13]));
    end
  endgenerate

  ////ROW 014
  generate
    localparam integer j14 = 14;
    for (i14 = 0; i14 < 24; i14 = i14 + 1)
    begin: addbit14
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j14+0][i14+0]), .Out(multi14[0][i14]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j14+0][i14+1]), .Out(multi14[1][i14]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j14+0][i14+2]), .Out(multi14[2][i14]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j14+0][i14+3]), .Out(multi14[3][i14]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j14+0][i14+4]), .Out(multi14[4][i14]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j14+1][i14+0]), .Out(multi14[5][i14]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j14+1][i14+1]), .Out(multi14[6][i14]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j14+1][i14+2]), .Out(multi14[7][i14]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j14+1][i14+3]), .Out(multi14[8][i14]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j14+1][i14+4]), .Out(multi14[9][i14]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j14+2][i14+0]), .Out(multi14[10][i14]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j14+2][i14+1]), .Out(multi14[11][i14]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j14+2][i14+2]), .Out(multi14[12][i14]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j14+2][i14+3]), .Out(multi14[13][i14]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j14+2][i14+4]), .Out(multi14[14][i14]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j14+3][i14+0]), .Out(multi14[15][i14]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j14+3][i14+1]), .Out(multi14[16][i14]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j14+3][i14+2]), .Out(multi14[17][i14]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j14+3][i14+3]), .Out(multi14[18][i14]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j14+3][i14+4]), .Out(multi14[19][i14]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j14+4][i14+0]), .Out(multi14[20][i14]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j14+4][i14+1]), .Out(multi14[21][i14]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j14+4][i14+2]), .Out(multi14[22][i14]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j14+4][i14+3]), .Out(multi14[23][i14]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j14+4][i14+4]), .Out(multi14[24][i14]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi14[0][i14]), .B(multi14[1][i14]), .Out(sum14[0][i14]));
      FP16_Add stage026(.A(multi14[2][i14]), .B(multi14[3][i14]), .Out(sum14[1][i14]));
      FP16_Add stage027(.A(multi14[4][i14]), .B(multi14[5][i14]), .Out(sum14[2][i14]));
      FP16_Add stage028(.A(multi14[6][i14]), .B(multi14[7][i14]), .Out(sum14[3][i14]));
      FP16_Add stage029(.A(multi14[8][i14]), .B(multi14[9][i14]), .Out(sum14[4][i14]));
      FP16_Add stage030(.A(multi14[10][i14]), .B(multi14[11][i14]), .Out(sum14[5][i14]));
      FP16_Add stage031(.A(multi14[12][i14]), .B(multi14[13][i14]), .Out(sum14[6][i14]));
      FP16_Add stage032(.A(multi14[14][i14]), .B(multi14[15][i14]), .Out(sum14[7][i14]));
      FP16_Add stage033(.A(multi14[16][i14]), .B(multi14[17][i14]), .Out(sum14[8][i14]));
      FP16_Add stage034(.A(multi14[18][i14]), .B(multi14[19][i14]), .Out(sum14[9][i14]));
      FP16_Add stage035(.A(multi14[20][i14]), .B(multi14[21][i14]), .Out(sum14[10][i14]));
      FP16_Add stage036(.A(multi14[22][i14]), .B(multi14[23][i14]), .Out(sum14[11][i14]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum14[0][i14]), .B(sum14[1][i14]), .Out(sum14[12][i14]));
      FP16_Add stage038(.A(sum14[2][i14]), .B(sum14[3][i14]), .Out(sum14[13][i14]));
      FP16_Add stage039(.A(sum14[4][i14]), .B(sum14[5][i14]), .Out(sum14[14][i14]));
      FP16_Add stage040(.A(sum14[6][i14]), .B(sum14[7][i14]), .Out(sum14[15][i14]));
      FP16_Add stage041(.A(sum14[8][i14]), .B(sum14[9][i14]), .Out(sum14[16][i14]));
      FP16_Add stage042(.A(sum14[10][i14]), .B(sum14[11][i14]), .Out(sum14[17][i14]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum14[12][i14]), .B(sum14[13][i14]), .Out(sum14[18][i14]));
      FP16_Add stage044(.A(sum14[14][i14]), .B(sum14[15][i14]), .Out(sum14[19][i14]));
      FP16_Add stage045(.A(sum14[16][i14]), .B(sum14[17][i14]), .Out(sum14[20][i14]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum14[18][i14]), .B(sum14[19][i14]), .Out(sum14[21][i14]));
      FP16_Add stage047(.A(sum14[20][i14]), .B(multi14[24][i14]), .Out(sum14[22][i14]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum14[21][i14]), .B(sum14[22][i14]), .Out(sum14[23][i14]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum14[23][i14]), .B(feature4Bias), .Out(data_11_array[j14][i14]));
    end
  endgenerate

  ////ROW 15
  generate
    localparam integer j15 = 15;
    for (i15 = 0; i15 < 24; i15 = i15 + 1)
    begin: addbit15
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j15+0][i15+0]), .Out(multi15[0][i15]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j15+0][i15+1]), .Out(multi15[1][i15]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j15+0][i15+2]), .Out(multi15[2][i15]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j15+0][i15+3]), .Out(multi15[3][i15]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j15+0][i15+4]), .Out(multi15[4][i15]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j15+1][i15+0]), .Out(multi15[5][i15]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j15+1][i15+1]), .Out(multi15[6][i15]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j15+1][i15+2]), .Out(multi15[7][i15]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j15+1][i15+3]), .Out(multi15[8][i15]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j15+1][i15+4]), .Out(multi15[9][i15]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j15+2][i15+0]), .Out(multi15[10][i15]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j15+2][i15+1]), .Out(multi15[11][i15]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j15+2][i15+2]), .Out(multi15[12][i15]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j15+2][i15+3]), .Out(multi15[13][i15]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j15+2][i15+4]), .Out(multi15[14][i15]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j15+3][i15+0]), .Out(multi15[15][i15]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j15+3][i15+1]), .Out(multi15[16][i15]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j15+3][i15+2]), .Out(multi15[17][i15]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j15+3][i15+3]), .Out(multi15[18][i15]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j15+3][i15+4]), .Out(multi15[19][i15]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j15+4][i15+0]), .Out(multi15[20][i15]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j15+4][i15+1]), .Out(multi15[21][i15]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j15+4][i15+2]), .Out(multi15[22][i15]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j15+4][i15+3]), .Out(multi15[23][i15]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j15+4][i15+4]), .Out(multi15[24][i15]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi15[0][i15]), .B(multi15[1][i15]), .Out(sum15[0][i15]));
      FP16_Add stage026(.A(multi15[2][i15]), .B(multi15[3][i15]), .Out(sum15[1][i15]));
      FP16_Add stage027(.A(multi15[4][i15]), .B(multi15[5][i15]), .Out(sum15[2][i15]));
      FP16_Add stage028(.A(multi15[6][i15]), .B(multi15[7][i15]), .Out(sum15[3][i15]));
      FP16_Add stage029(.A(multi15[8][i15]), .B(multi15[9][i15]), .Out(sum15[4][i15]));
      FP16_Add stage030(.A(multi15[10][i15]), .B(multi15[11][i15]), .Out(sum15[5][i15]));
      FP16_Add stage031(.A(multi15[12][i15]), .B(multi15[13][i15]), .Out(sum15[6][i15]));
      FP16_Add stage032(.A(multi15[14][i15]), .B(multi15[15][i15]), .Out(sum15[7][i15]));
      FP16_Add stage033(.A(multi15[16][i15]), .B(multi15[17][i15]), .Out(sum15[8][i15]));
      FP16_Add stage034(.A(multi15[18][i15]), .B(multi15[19][i15]), .Out(sum15[9][i15]));
      FP16_Add stage035(.A(multi15[20][i15]), .B(multi15[21][i15]), .Out(sum15[10][i15]));
      FP16_Add stage036(.A(multi15[22][i15]), .B(multi15[23][i15]), .Out(sum15[11][i15]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum15[0][i15]), .B(sum15[1][i15]), .Out(sum15[12][i15]));
      FP16_Add stage038(.A(sum15[2][i15]), .B(sum15[3][i15]), .Out(sum15[13][i15]));
      FP16_Add stage039(.A(sum15[4][i15]), .B(sum15[5][i15]), .Out(sum15[14][i15]));
      FP16_Add stage040(.A(sum15[6][i15]), .B(sum15[7][i15]), .Out(sum15[15][i15]));
      FP16_Add stage041(.A(sum15[8][i15]), .B(sum15[9][i15]), .Out(sum15[16][i15]));
      FP16_Add stage042(.A(sum15[10][i15]), .B(sum15[11][i15]), .Out(sum15[17][i15]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum15[12][i15]), .B(sum15[13][i15]), .Out(sum15[18][i15]));
      FP16_Add stage044(.A(sum15[14][i15]), .B(sum15[15][i15]), .Out(sum15[19][i15]));
      FP16_Add stage045(.A(sum15[16][i15]), .B(sum15[17][i15]), .Out(sum15[20][i15]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum15[18][i15]), .B(sum15[19][i15]), .Out(sum15[21][i15]));
      FP16_Add stage047(.A(sum15[20][i15]), .B(multi15[24][i15]), .Out(sum15[22][i15]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum15[21][i15]), .B(sum15[22][i15]), .Out(sum15[23][i15]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum15[23][i15]), .B(feature4Bias), .Out(data_11_array[j15][i15]));
    end
  endgenerate
  
  ////ROW 16
  generate
    localparam integer j16 = 16;
    for (i16 = 0; i16 < 24; i16 = i16 + 1)
    begin: addbit16
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j16+0][i16+0]), .Out(multi16[0][i16]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j16+0][i16+1]), .Out(multi16[1][i16]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j16+0][i16+2]), .Out(multi16[2][i16]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j16+0][i16+3]), .Out(multi16[3][i16]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j16+0][i16+4]), .Out(multi16[4][i16]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j16+1][i16+0]), .Out(multi16[5][i16]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j16+1][i16+1]), .Out(multi16[6][i16]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j16+1][i16+2]), .Out(multi16[7][i16]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j16+1][i16+3]), .Out(multi16[8][i16]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j16+1][i16+4]), .Out(multi16[9][i16]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j16+2][i16+0]), .Out(multi16[10][i16]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j16+2][i16+1]), .Out(multi16[11][i16]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j16+2][i16+2]), .Out(multi16[12][i16]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j16+2][i16+3]), .Out(multi16[13][i16]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j16+2][i16+4]), .Out(multi16[14][i16]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j16+3][i16+0]), .Out(multi16[15][i16]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j16+3][i16+1]), .Out(multi16[16][i16]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j16+3][i16+2]), .Out(multi16[17][i16]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j16+3][i16+3]), .Out(multi16[18][i16]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j16+3][i16+4]), .Out(multi16[19][i16]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j16+4][i16+0]), .Out(multi16[20][i16]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j16+4][i16+1]), .Out(multi16[21][i16]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j16+4][i16+2]), .Out(multi16[22][i16]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j16+4][i16+3]), .Out(multi16[23][i16]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j16+4][i16+4]), .Out(multi16[24][i16]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi16[0][i16]), .B(multi16[1][i16]), .Out(sum16[0][i16]));
      FP16_Add stage026(.A(multi16[2][i16]), .B(multi16[3][i16]), .Out(sum16[1][i16]));
      FP16_Add stage027(.A(multi16[4][i16]), .B(multi16[5][i16]), .Out(sum16[2][i16]));
      FP16_Add stage028(.A(multi16[6][i16]), .B(multi16[7][i16]), .Out(sum16[3][i16]));
      FP16_Add stage029(.A(multi16[8][i16]), .B(multi16[9][i16]), .Out(sum16[4][i16]));
      FP16_Add stage030(.A(multi16[10][i16]), .B(multi16[11][i16]), .Out(sum16[5][i16]));
      FP16_Add stage031(.A(multi16[12][i16]), .B(multi16[13][i16]), .Out(sum16[6][i16]));
      FP16_Add stage032(.A(multi16[14][i16]), .B(multi16[15][i16]), .Out(sum16[7][i16]));
      FP16_Add stage033(.A(multi16[16][i16]), .B(multi16[17][i16]), .Out(sum16[8][i16]));
      FP16_Add stage034(.A(multi16[18][i16]), .B(multi16[19][i16]), .Out(sum16[9][i16]));
      FP16_Add stage035(.A(multi16[20][i16]), .B(multi16[21][i16]), .Out(sum16[10][i16]));
      FP16_Add stage036(.A(multi16[22][i16]), .B(multi16[23][i16]), .Out(sum16[11][i16]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum16[0][i16]), .B(sum16[1][i16]), .Out(sum16[12][i16]));
      FP16_Add stage038(.A(sum16[2][i16]), .B(sum16[3][i16]), .Out(sum16[13][i16]));
      FP16_Add stage039(.A(sum16[4][i16]), .B(sum16[5][i16]), .Out(sum16[14][i16]));
      FP16_Add stage040(.A(sum16[6][i16]), .B(sum16[7][i16]), .Out(sum16[15][i16]));
      FP16_Add stage041(.A(sum16[8][i16]), .B(sum16[9][i16]), .Out(sum16[16][i16]));
      FP16_Add stage042(.A(sum16[10][i16]), .B(sum16[11][i16]), .Out(sum16[17][i16]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum16[12][i16]), .B(sum16[13][i16]), .Out(sum16[18][i16]));
      FP16_Add stage044(.A(sum16[14][i16]), .B(sum16[15][i16]), .Out(sum16[19][i16]));
      FP16_Add stage045(.A(sum16[16][i16]), .B(sum16[17][i16]), .Out(sum16[20][i16]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum16[18][i16]), .B(sum16[19][i16]), .Out(sum16[21][i16]));
      FP16_Add stage047(.A(sum16[20][i16]), .B(multi16[24][i16]), .Out(sum16[22][i16]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum16[21][i16]), .B(sum16[22][i16]), .Out(sum16[23][i16]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum16[23][i16]), .B(feature4Bias), .Out(data_11_array[j16][i16]));
    end
  endgenerate
  
  ////ROW 17
  generate
    localparam integer j17 = 17;
    for (i17 = 0; i17 < 24; i17 = i17 + 1)
    begin: addbit17
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j17+0][i17+0]), .Out(multi17[0][i17]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j17+0][i17+1]), .Out(multi17[1][i17]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j17+0][i17+2]), .Out(multi17[2][i17]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j17+0][i17+3]), .Out(multi17[3][i17]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j17+0][i17+4]), .Out(multi17[4][i17]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j17+1][i17+0]), .Out(multi17[5][i17]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j17+1][i17+1]), .Out(multi17[6][i17]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j17+1][i17+2]), .Out(multi17[7][i17]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j17+1][i17+3]), .Out(multi17[8][i17]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j17+1][i17+4]), .Out(multi17[9][i17]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j17+2][i17+0]), .Out(multi17[10][i17]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j17+2][i17+1]), .Out(multi17[11][i17]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j17+2][i17+2]), .Out(multi17[12][i17]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j17+2][i17+3]), .Out(multi17[13][i17]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j17+2][i17+4]), .Out(multi17[14][i17]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j17+3][i17+0]), .Out(multi17[15][i17]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j17+3][i17+1]), .Out(multi17[16][i17]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j17+3][i17+2]), .Out(multi17[17][i17]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j17+3][i17+3]), .Out(multi17[18][i17]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j17+3][i17+4]), .Out(multi17[19][i17]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j17+4][i17+0]), .Out(multi17[20][i17]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j17+4][i17+1]), .Out(multi17[21][i17]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j17+4][i17+2]), .Out(multi17[22][i17]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j17+4][i17+3]), .Out(multi17[23][i17]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j17+4][i17+4]), .Out(multi17[24][i17]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi17[0][i17]), .B(multi17[1][i17]), .Out(sum17[0][i17]));
      FP16_Add stage026(.A(multi17[2][i17]), .B(multi17[3][i17]), .Out(sum17[1][i17]));
      FP16_Add stage027(.A(multi17[4][i17]), .B(multi17[5][i17]), .Out(sum17[2][i17]));
      FP16_Add stage028(.A(multi17[6][i17]), .B(multi17[7][i17]), .Out(sum17[3][i17]));
      FP16_Add stage029(.A(multi17[8][i17]), .B(multi17[9][i17]), .Out(sum17[4][i17]));
      FP16_Add stage030(.A(multi17[10][i17]), .B(multi17[11][i17]), .Out(sum17[5][i17]));
      FP16_Add stage031(.A(multi17[12][i17]), .B(multi17[13][i17]), .Out(sum17[6][i17]));
      FP16_Add stage032(.A(multi17[14][i17]), .B(multi17[15][i17]), .Out(sum17[7][i17]));
      FP16_Add stage033(.A(multi17[16][i17]), .B(multi17[17][i17]), .Out(sum17[8][i17]));
      FP16_Add stage034(.A(multi17[18][i17]), .B(multi17[19][i17]), .Out(sum17[9][i17]));
      FP16_Add stage035(.A(multi17[20][i17]), .B(multi17[21][i17]), .Out(sum17[10][i17]));
      FP16_Add stage036(.A(multi17[22][i17]), .B(multi17[23][i17]), .Out(sum17[11][i17]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum17[0][i17]), .B(sum17[1][i17]), .Out(sum17[12][i17]));
      FP16_Add stage038(.A(sum17[2][i17]), .B(sum17[3][i17]), .Out(sum17[13][i17]));
      FP16_Add stage039(.A(sum17[4][i17]), .B(sum17[5][i17]), .Out(sum17[14][i17]));
      FP16_Add stage040(.A(sum17[6][i17]), .B(sum17[7][i17]), .Out(sum17[15][i17]));
      FP16_Add stage041(.A(sum17[8][i17]), .B(sum17[9][i17]), .Out(sum17[16][i17]));
      FP16_Add stage042(.A(sum17[10][i17]), .B(sum17[11][i17]), .Out(sum17[17][i17]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum17[12][i17]), .B(sum17[13][i17]), .Out(sum17[18][i17]));
      FP16_Add stage044(.A(sum17[14][i17]), .B(sum17[15][i17]), .Out(sum17[19][i17]));
      FP16_Add stage045(.A(sum17[16][i17]), .B(sum17[17][i17]), .Out(sum17[20][i17]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum17[18][i17]), .B(sum17[19][i17]), .Out(sum17[21][i17]));
      FP16_Add stage047(.A(sum17[20][i17]), .B(multi17[24][i17]), .Out(sum17[22][i17]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum17[21][i17]), .B(sum17[22][i17]), .Out(sum17[23][i17]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum17[23][i17]), .B(feature4Bias), .Out(data_11_array[j17][i17]));
    end
  endgenerate

////ROW 18
  generate
    localparam integer j18 = 18;
    for (i18 = 0; i18 < 24; i18 = i18 + 1)
    begin: addbit18
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j18+0][i18+0]), .Out(multi18[0][i18]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j18+0][i18+1]), .Out(multi18[1][i18]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j18+0][i18+2]), .Out(multi18[2][i18]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j18+0][i18+3]), .Out(multi18[3][i18]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j18+0][i18+4]), .Out(multi18[4][i18]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j18+1][i18+0]), .Out(multi18[5][i18]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j18+1][i18+1]), .Out(multi18[6][i18]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j18+1][i18+2]), .Out(multi18[7][i18]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j18+1][i18+3]), .Out(multi18[8][i18]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j18+1][i18+4]), .Out(multi18[9][i18]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j18+2][i18+0]), .Out(multi18[10][i18]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j18+2][i18+1]), .Out(multi18[11][i18]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j18+2][i18+2]), .Out(multi18[12][i18]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j18+2][i18+3]), .Out(multi18[13][i18]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j18+2][i18+4]), .Out(multi18[14][i18]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j18+3][i18+0]), .Out(multi18[15][i18]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j18+3][i18+1]), .Out(multi18[16][i18]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j18+3][i18+2]), .Out(multi18[17][i18]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j18+3][i18+3]), .Out(multi18[18][i18]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j18+3][i18+4]), .Out(multi18[19][i18]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j18+4][i18+0]), .Out(multi18[20][i18]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j18+4][i18+1]), .Out(multi18[21][i18]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j18+4][i18+2]), .Out(multi18[22][i18]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j18+4][i18+3]), .Out(multi18[23][i18]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j18+4][i18+4]), .Out(multi18[24][i18]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi18[0][i18]), .B(multi18[1][i18]), .Out(sum18[0][i18]));
      FP16_Add stage026(.A(multi18[2][i18]), .B(multi18[3][i18]), .Out(sum18[1][i18]));
      FP16_Add stage027(.A(multi18[4][i18]), .B(multi18[5][i18]), .Out(sum18[2][i18]));
      FP16_Add stage028(.A(multi18[6][i18]), .B(multi18[7][i18]), .Out(sum18[3][i18]));
      FP16_Add stage029(.A(multi18[8][i18]), .B(multi18[9][i18]), .Out(sum18[4][i18]));
      FP16_Add stage030(.A(multi18[10][i18]), .B(multi18[11][i18]), .Out(sum18[5][i18]));
      FP16_Add stage031(.A(multi18[12][i18]), .B(multi18[13][i18]), .Out(sum18[6][i18]));
      FP16_Add stage032(.A(multi18[14][i18]), .B(multi18[15][i18]), .Out(sum18[7][i18]));
      FP16_Add stage033(.A(multi18[16][i18]), .B(multi18[17][i18]), .Out(sum18[8][i18]));
      FP16_Add stage034(.A(multi18[18][i18]), .B(multi18[19][i18]), .Out(sum18[9][i18]));
      FP16_Add stage035(.A(multi18[20][i18]), .B(multi18[21][i18]), .Out(sum18[10][i18]));
      FP16_Add stage036(.A(multi18[22][i18]), .B(multi18[23][i18]), .Out(sum18[11][i18]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum18[0][i18]), .B(sum18[1][i18]), .Out(sum18[12][i18]));
      FP16_Add stage038(.A(sum18[2][i18]), .B(sum18[3][i18]), .Out(sum18[13][i18]));
      FP16_Add stage039(.A(sum18[4][i18]), .B(sum18[5][i18]), .Out(sum18[14][i18]));
      FP16_Add stage040(.A(sum18[6][i18]), .B(sum18[7][i18]), .Out(sum18[15][i18]));
      FP16_Add stage041(.A(sum18[8][i18]), .B(sum18[9][i18]), .Out(sum18[16][i18]));
      FP16_Add stage042(.A(sum18[10][i18]), .B(sum18[11][i18]), .Out(sum18[17][i18]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum18[12][i18]), .B(sum18[13][i18]), .Out(sum18[18][i18]));
      FP16_Add stage044(.A(sum18[14][i18]), .B(sum18[15][i18]), .Out(sum18[19][i18]));
      FP16_Add stage045(.A(sum18[16][i18]), .B(sum18[17][i18]), .Out(sum18[20][i18]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum18[18][i18]), .B(sum18[19][i18]), .Out(sum18[21][i18]));
      FP16_Add stage047(.A(sum18[20][i18]), .B(multi18[24][i18]), .Out(sum18[22][i18]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum18[21][i18]), .B(sum18[22][i18]), .Out(sum18[23][i18]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum18[23][i18]), .B(feature4Bias), .Out(data_11_array[j18][i18]));
    end
  endgenerate

////ROW 19
  generate
    localparam integer j19 = 19;
    for (i19 = 0; i19 < 24; i19 = i19 + 1)
    begin: addbit19
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j19+0][i19+0]), .Out(multi19[0][i19]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j19+0][i19+1]), .Out(multi19[1][i19]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j19+0][i19+2]), .Out(multi19[2][i19]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j19+0][i19+3]), .Out(multi19[3][i19]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j19+0][i19+4]), .Out(multi19[4][i19]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j19+1][i19+0]), .Out(multi19[5][i19]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j19+1][i19+1]), .Out(multi19[6][i19]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j19+1][i19+2]), .Out(multi19[7][i19]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j19+1][i19+3]), .Out(multi19[8][i19]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j19+1][i19+4]), .Out(multi19[9][i19]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j19+2][i19+0]), .Out(multi19[10][i19]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j19+2][i19+1]), .Out(multi19[11][i19]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j19+2][i19+2]), .Out(multi19[12][i19]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j19+2][i19+3]), .Out(multi19[13][i19]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j19+2][i19+4]), .Out(multi19[14][i19]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j19+3][i19+0]), .Out(multi19[15][i19]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j19+3][i19+1]), .Out(multi19[16][i19]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j19+3][i19+2]), .Out(multi19[17][i19]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j19+3][i19+3]), .Out(multi19[18][i19]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j19+3][i19+4]), .Out(multi19[19][i19]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j19+4][i19+0]), .Out(multi19[20][i19]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j19+4][i19+1]), .Out(multi19[21][i19]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j19+4][i19+2]), .Out(multi19[22][i19]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j19+4][i19+3]), .Out(multi19[23][i19]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j19+4][i19+4]), .Out(multi19[24][i19]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi19[0][i19]), .B(multi19[1][i19]), .Out(sum19[0][i19]));
      FP16_Add stage026(.A(multi19[2][i19]), .B(multi19[3][i19]), .Out(sum19[1][i19]));
      FP16_Add stage027(.A(multi19[4][i19]), .B(multi19[5][i19]), .Out(sum19[2][i19]));
      FP16_Add stage028(.A(multi19[6][i19]), .B(multi19[7][i19]), .Out(sum19[3][i19]));
      FP16_Add stage029(.A(multi19[8][i19]), .B(multi19[9][i19]), .Out(sum19[4][i19]));
      FP16_Add stage030(.A(multi19[10][i19]), .B(multi19[11][i19]), .Out(sum19[5][i19]));
      FP16_Add stage031(.A(multi19[12][i19]), .B(multi19[13][i19]), .Out(sum19[6][i19]));
      FP16_Add stage032(.A(multi19[14][i19]), .B(multi19[15][i19]), .Out(sum19[7][i19]));
      FP16_Add stage033(.A(multi19[16][i19]), .B(multi19[17][i19]), .Out(sum19[8][i19]));
      FP16_Add stage034(.A(multi19[18][i19]), .B(multi19[19][i19]), .Out(sum19[9][i19]));
      FP16_Add stage035(.A(multi19[20][i19]), .B(multi19[21][i19]), .Out(sum19[10][i19]));
      FP16_Add stage036(.A(multi19[22][i19]), .B(multi19[23][i19]), .Out(sum19[11][i19]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum19[0][i19]), .B(sum19[1][i19]), .Out(sum19[12][i19]));
      FP16_Add stage038(.A(sum19[2][i19]), .B(sum19[3][i19]), .Out(sum19[13][i19]));
      FP16_Add stage039(.A(sum19[4][i19]), .B(sum19[5][i19]), .Out(sum19[14][i19]));
      FP16_Add stage040(.A(sum19[6][i19]), .B(sum19[7][i19]), .Out(sum19[15][i19]));
      FP16_Add stage041(.A(sum19[8][i19]), .B(sum19[9][i19]), .Out(sum19[16][i19]));
      FP16_Add stage042(.A(sum19[10][i19]), .B(sum19[11][i19]), .Out(sum19[17][i19]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum19[12][i19]), .B(sum19[13][i19]), .Out(sum19[18][i19]));
      FP16_Add stage044(.A(sum19[14][i19]), .B(sum19[15][i19]), .Out(sum19[19][i19]));
      FP16_Add stage045(.A(sum19[16][i19]), .B(sum19[17][i19]), .Out(sum19[20][i19]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum19[18][i19]), .B(sum19[19][i19]), .Out(sum19[21][i19]));
      FP16_Add stage047(.A(sum19[20][i19]), .B(multi19[24][i19]), .Out(sum19[22][i19]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum19[21][i19]), .B(sum19[22][i19]), .Out(sum19[23][i19]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum19[23][i19]), .B(feature4Bias), .Out(data_11_array[j19][i19]));
    end
  endgenerate

////ROW 20
  generate
    localparam integer j20 = 20;
    for (i20 = 0; i20 < 24; i20 = i20 + 1)
    begin: addbit20
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j20+0][i20+0]), .Out(multi20[0][i20]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j20+0][i20+1]), .Out(multi20[1][i20]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j20+0][i20+2]), .Out(multi20[2][i20]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j20+0][i20+3]), .Out(multi20[3][i20]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j20+0][i20+4]), .Out(multi20[4][i20]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j20+1][i20+0]), .Out(multi20[5][i20]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j20+1][i20+1]), .Out(multi20[6][i20]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j20+1][i20+2]), .Out(multi20[7][i20]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j20+1][i20+3]), .Out(multi20[8][i20]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j20+1][i20+4]), .Out(multi20[9][i20]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j20+2][i20+0]), .Out(multi20[10][i20]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j20+2][i20+1]), .Out(multi20[11][i20]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j20+2][i20+2]), .Out(multi20[12][i20]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j20+2][i20+3]), .Out(multi20[13][i20]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j20+2][i20+4]), .Out(multi20[14][i20]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j20+3][i20+0]), .Out(multi20[15][i20]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j20+3][i20+1]), .Out(multi20[16][i20]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j20+3][i20+2]), .Out(multi20[17][i20]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j20+3][i20+3]), .Out(multi20[18][i20]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j20+3][i20+4]), .Out(multi20[19][i20]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j20+4][i20+0]), .Out(multi20[20][i20]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j20+4][i20+1]), .Out(multi20[21][i20]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j20+4][i20+2]), .Out(multi20[22][i20]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j20+4][i20+3]), .Out(multi20[23][i20]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j20+4][i20+4]), .Out(multi20[24][i20]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi20[0][i20]), .B(multi20[1][i20]), .Out(sum20[0][i20]));
      FP16_Add stage026(.A(multi20[2][i20]), .B(multi20[3][i20]), .Out(sum20[1][i20]));
      FP16_Add stage027(.A(multi20[4][i20]), .B(multi20[5][i20]), .Out(sum20[2][i20]));
      FP16_Add stage028(.A(multi20[6][i20]), .B(multi20[7][i20]), .Out(sum20[3][i20]));
      FP16_Add stage029(.A(multi20[8][i20]), .B(multi20[9][i20]), .Out(sum20[4][i20]));
      FP16_Add stage030(.A(multi20[10][i20]), .B(multi20[11][i20]), .Out(sum20[5][i20]));
      FP16_Add stage031(.A(multi20[12][i20]), .B(multi20[13][i20]), .Out(sum20[6][i20]));
      FP16_Add stage032(.A(multi20[14][i20]), .B(multi20[15][i20]), .Out(sum20[7][i20]));
      FP16_Add stage033(.A(multi20[16][i20]), .B(multi20[17][i20]), .Out(sum20[8][i20]));
      FP16_Add stage034(.A(multi20[18][i20]), .B(multi20[19][i20]), .Out(sum20[9][i20]));
      FP16_Add stage035(.A(multi20[20][i20]), .B(multi20[21][i20]), .Out(sum20[10][i20]));
      FP16_Add stage036(.A(multi20[22][i20]), .B(multi20[23][i20]), .Out(sum20[11][i20]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum20[0][i20]), .B(sum20[1][i20]), .Out(sum20[12][i20]));
      FP16_Add stage038(.A(sum20[2][i20]), .B(sum20[3][i20]), .Out(sum20[13][i20]));
      FP16_Add stage039(.A(sum20[4][i20]), .B(sum20[5][i20]), .Out(sum20[14][i20]));
      FP16_Add stage040(.A(sum20[6][i20]), .B(sum20[7][i20]), .Out(sum20[15][i20]));
      FP16_Add stage041(.A(sum20[8][i20]), .B(sum20[9][i20]), .Out(sum20[16][i20]));
      FP16_Add stage042(.A(sum20[10][i20]), .B(sum20[11][i20]), .Out(sum20[17][i20]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum20[12][i20]), .B(sum20[13][i20]), .Out(sum20[18][i20]));
      FP16_Add stage044(.A(sum20[14][i20]), .B(sum20[15][i20]), .Out(sum20[19][i20]));
      FP16_Add stage045(.A(sum20[16][i20]), .B(sum20[17][i20]), .Out(sum20[20][i20]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum20[18][i20]), .B(sum20[19][i20]), .Out(sum20[21][i20]));
      FP16_Add stage047(.A(sum20[20][i20]), .B(multi20[24][i20]), .Out(sum20[22][i20]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum20[21][i20]), .B(sum20[22][i20]), .Out(sum20[23][i20]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum20[23][i20]), .B(feature4Bias), .Out(data_11_array[j20][i20]));
    end
  endgenerate

////ROW 21
  generate
    localparam integer j21 = 21;
    for (i21 = 0; i21 < 24; i21 = i21 + 1)
    begin: addbit21
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j21+0][i21+0]), .Out(multi21[0][i21]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j21+0][i21+1]), .Out(multi21[1][i21]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j21+0][i21+2]), .Out(multi21[2][i21]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j21+0][i21+3]), .Out(multi21[3][i21]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j21+0][i21+4]), .Out(multi21[4][i21]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j21+1][i21+0]), .Out(multi21[5][i21]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j21+1][i21+1]), .Out(multi21[6][i21]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j21+1][i21+2]), .Out(multi21[7][i21]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j21+1][i21+3]), .Out(multi21[8][i21]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j21+1][i21+4]), .Out(multi21[9][i21]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j21+2][i21+0]), .Out(multi21[10][i21]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j21+2][i21+1]), .Out(multi21[11][i21]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j21+2][i21+2]), .Out(multi21[12][i21]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j21+2][i21+3]), .Out(multi21[13][i21]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j21+2][i21+4]), .Out(multi21[14][i21]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j21+3][i21+0]), .Out(multi21[15][i21]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j21+3][i21+1]), .Out(multi21[16][i21]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j21+3][i21+2]), .Out(multi21[17][i21]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j21+3][i21+3]), .Out(multi21[18][i21]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j21+3][i21+4]), .Out(multi21[19][i21]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j21+4][i21+0]), .Out(multi21[20][i21]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j21+4][i21+1]), .Out(multi21[21][i21]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j21+4][i21+2]), .Out(multi21[22][i21]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j21+4][i21+3]), .Out(multi21[23][i21]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j21+4][i21+4]), .Out(multi21[24][i21]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi21[0][i21]), .B(multi21[1][i21]), .Out(sum21[0][i21]));
      FP16_Add stage026(.A(multi21[2][i21]), .B(multi21[3][i21]), .Out(sum21[1][i21]));
      FP16_Add stage027(.A(multi21[4][i21]), .B(multi21[5][i21]), .Out(sum21[2][i21]));
      FP16_Add stage028(.A(multi21[6][i21]), .B(multi21[7][i21]), .Out(sum21[3][i21]));
      FP16_Add stage029(.A(multi21[8][i21]), .B(multi21[9][i21]), .Out(sum21[4][i21]));
      FP16_Add stage030(.A(multi21[10][i21]), .B(multi21[11][i21]), .Out(sum21[5][i21]));
      FP16_Add stage031(.A(multi21[12][i21]), .B(multi21[13][i21]), .Out(sum21[6][i21]));
      FP16_Add stage032(.A(multi21[14][i21]), .B(multi21[15][i21]), .Out(sum21[7][i21]));
      FP16_Add stage033(.A(multi21[16][i21]), .B(multi21[17][i21]), .Out(sum21[8][i21]));
      FP16_Add stage034(.A(multi21[18][i21]), .B(multi21[19][i21]), .Out(sum21[9][i21]));
      FP16_Add stage035(.A(multi21[20][i21]), .B(multi21[21][i21]), .Out(sum21[10][i21]));
      FP16_Add stage036(.A(multi21[22][i21]), .B(multi21[23][i21]), .Out(sum21[11][i21]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum21[0][i21]), .B(sum21[1][i21]), .Out(sum21[12][i21]));
      FP16_Add stage038(.A(sum21[2][i21]), .B(sum21[3][i21]), .Out(sum21[13][i21]));
      FP16_Add stage039(.A(sum21[4][i21]), .B(sum21[5][i21]), .Out(sum21[14][i21]));
      FP16_Add stage040(.A(sum21[6][i21]), .B(sum21[7][i21]), .Out(sum21[15][i21]));
      FP16_Add stage041(.A(sum21[8][i21]), .B(sum21[9][i21]), .Out(sum21[16][i21]));
      FP16_Add stage042(.A(sum21[10][i21]), .B(sum21[11][i21]), .Out(sum21[17][i21]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum21[12][i21]), .B(sum21[13][i21]), .Out(sum21[18][i21]));
      FP16_Add stage044(.A(sum21[14][i21]), .B(sum21[15][i21]), .Out(sum21[19][i21]));
      FP16_Add stage045(.A(sum21[16][i21]), .B(sum21[17][i21]), .Out(sum21[20][i21]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum21[18][i21]), .B(sum21[19][i21]), .Out(sum21[21][i21]));
      FP16_Add stage047(.A(sum21[20][i21]), .B(multi21[24][i21]), .Out(sum21[22][i21]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum21[21][i21]), .B(sum21[22][i21]), .Out(sum21[23][i21]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum21[23][i21]), .B(feature4Bias), .Out(data_11_array[j21][i21]));
    end
  endgenerate

////ROW 22
  generate
    localparam integer j22 = 22;
    for (i22 = 0; i22 < 24; i22 = i22 + 1)
    begin: addbit22
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j22+0][i22+0]), .Out(multi22[0][i22]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j22+0][i22+1]), .Out(multi22[1][i22]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j22+0][i22+2]), .Out(multi22[2][i22]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j22+0][i22+3]), .Out(multi22[3][i22]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j22+0][i22+4]), .Out(multi22[4][i22]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j22+1][i22+0]), .Out(multi22[5][i22]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j22+1][i22+1]), .Out(multi22[6][i22]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j22+1][i22+2]), .Out(multi22[7][i22]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j22+1][i22+3]), .Out(multi22[8][i22]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j22+1][i22+4]), .Out(multi22[9][i22]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j22+2][i22+0]), .Out(multi22[10][i22]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j22+2][i22+1]), .Out(multi22[11][i22]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j22+2][i22+2]), .Out(multi22[12][i22]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j22+2][i22+3]), .Out(multi22[13][i22]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j22+2][i22+4]), .Out(multi22[14][i22]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j22+3][i22+0]), .Out(multi22[15][i22]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j22+3][i22+1]), .Out(multi22[16][i22]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j22+3][i22+2]), .Out(multi22[17][i22]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j22+3][i22+3]), .Out(multi22[18][i22]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j22+3][i22+4]), .Out(multi22[19][i22]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j22+4][i22+0]), .Out(multi22[20][i22]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j22+4][i22+1]), .Out(multi22[21][i22]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j22+4][i22+2]), .Out(multi22[22][i22]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j22+4][i22+3]), .Out(multi22[23][i22]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j22+4][i22+4]), .Out(multi22[24][i22]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi22[0][i22]), .B(multi22[1][i22]), .Out(sum22[0][i22]));
      FP16_Add stage026(.A(multi22[2][i22]), .B(multi22[3][i22]), .Out(sum22[1][i22]));
      FP16_Add stage027(.A(multi22[4][i22]), .B(multi22[5][i22]), .Out(sum22[2][i22]));
      FP16_Add stage028(.A(multi22[6][i22]), .B(multi22[7][i22]), .Out(sum22[3][i22]));
      FP16_Add stage029(.A(multi22[8][i22]), .B(multi22[9][i22]), .Out(sum22[4][i22]));
      FP16_Add stage030(.A(multi22[10][i22]), .B(multi22[11][i22]), .Out(sum22[5][i22]));
      FP16_Add stage031(.A(multi22[12][i22]), .B(multi22[13][i22]), .Out(sum22[6][i22]));
      FP16_Add stage032(.A(multi22[14][i22]), .B(multi22[15][i22]), .Out(sum22[7][i22]));
      FP16_Add stage033(.A(multi22[16][i22]), .B(multi22[17][i22]), .Out(sum22[8][i22]));
      FP16_Add stage034(.A(multi22[18][i22]), .B(multi22[19][i22]), .Out(sum22[9][i22]));
      FP16_Add stage035(.A(multi22[20][i22]), .B(multi22[21][i22]), .Out(sum22[10][i22]));
      FP16_Add stage036(.A(multi22[22][i22]), .B(multi22[23][i22]), .Out(sum22[11][i22]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum22[0][i22]), .B(sum22[1][i22]), .Out(sum22[12][i22]));
      FP16_Add stage038(.A(sum22[2][i22]), .B(sum22[3][i22]), .Out(sum22[13][i22]));
      FP16_Add stage039(.A(sum22[4][i22]), .B(sum22[5][i22]), .Out(sum22[14][i22]));
      FP16_Add stage040(.A(sum22[6][i22]), .B(sum22[7][i22]), .Out(sum22[15][i22]));
      FP16_Add stage041(.A(sum22[8][i22]), .B(sum22[9][i22]), .Out(sum22[16][i22]));
      FP16_Add stage042(.A(sum22[10][i22]), .B(sum22[11][i22]), .Out(sum22[17][i22]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum22[12][i22]), .B(sum22[13][i22]), .Out(sum22[18][i22]));
      FP16_Add stage044(.A(sum22[14][i22]), .B(sum22[15][i22]), .Out(sum22[19][i22]));
      FP16_Add stage045(.A(sum22[16][i22]), .B(sum22[17][i22]), .Out(sum22[20][i22]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum22[18][i22]), .B(sum22[19][i22]), .Out(sum22[21][i22]));
      FP16_Add stage047(.A(sum22[20][i22]), .B(multi22[24][i22]), .Out(sum22[22][i22]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum22[21][i22]), .B(sum22[22][i22]), .Out(sum22[23][i22]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum22[23][i22]), .B(feature4Bias), .Out(data_11_array[j22][i22]));
    end
  endgenerate

////ROW 23
  generate
    localparam integer j23 = 23;
    for (i23 = 0; i23 < 24; i23 = i23 + 1)
    begin: addbit23
    
      ////Multiplication
      FP16_Multiply stage00(.A(feature4Weight_0), .B(data_array[j23+0][i23+0]), .Out(multi23[0][i23]));
      FP16_Multiply stage01(.A(feature4Weight_1), .B(data_array[j23+0][i23+1]), .Out(multi23[1][i23]));
      FP16_Multiply stage02(.A(feature4Weight_2), .B(data_array[j23+0][i23+2]), .Out(multi23[2][i23]));
      FP16_Multiply stage03(.A(feature4Weight_3), .B(data_array[j23+0][i23+3]), .Out(multi23[3][i23]));
      FP16_Multiply stage04(.A(feature4Weight_4), .B(data_array[j23+0][i23+4]), .Out(multi23[4][i23]));
      FP16_Multiply stage05(.A(feature4Weight_5), .B(data_array[j23+1][i23+0]), .Out(multi23[5][i23]));
      FP16_Multiply stage06(.A(feature4Weight_6), .B(data_array[j23+1][i23+1]), .Out(multi23[6][i23]));
      FP16_Multiply stage07(.A(feature4Weight_7), .B(data_array[j23+1][i23+2]), .Out(multi23[7][i23]));
      FP16_Multiply stage08(.A(feature4Weight_8), .B(data_array[j23+1][i23+3]), .Out(multi23[8][i23]));
      FP16_Multiply stage09(.A(feature4Weight_9), .B(data_array[j23+1][i23+4]), .Out(multi23[9][i23]));
      FP16_Multiply stage010(.A(feature4Weight_10), .B(data_array[j23+2][i23+0]), .Out(multi23[10][i23]));
      FP16_Multiply stage011(.A(feature4Weight_11), .B(data_array[j23+2][i23+1]), .Out(multi23[11][i23]));
      FP16_Multiply stage012(.A(feature4Weight_12), .B(data_array[j23+2][i23+2]), .Out(multi23[12][i23]));
      FP16_Multiply stage013(.A(feature4Weight_13), .B(data_array[j23+2][i23+3]), .Out(multi23[13][i23]));
      FP16_Multiply stage014(.A(feature4Weight_14), .B(data_array[j23+2][i23+4]), .Out(multi23[14][i23]));
      FP16_Multiply stage015(.A(feature4Weight_15), .B(data_array[j23+3][i23+0]), .Out(multi23[15][i23]));
      FP16_Multiply stage016(.A(feature4Weight_16), .B(data_array[j23+3][i23+1]), .Out(multi23[16][i23]));
      FP16_Multiply stage017(.A(feature4Weight_17), .B(data_array[j23+3][i23+2]), .Out(multi23[17][i23]));
      FP16_Multiply stage018(.A(feature4Weight_18), .B(data_array[j23+3][i23+3]), .Out(multi23[18][i23]));
      FP16_Multiply stage019(.A(feature4Weight_19), .B(data_array[j23+3][i23+4]), .Out(multi23[19][i23]));
      FP16_Multiply stage020(.A(feature4Weight_20), .B(data_array[j23+4][i23+0]), .Out(multi23[20][i23]));
      FP16_Multiply stage021(.A(feature4Weight_21), .B(data_array[j23+4][i23+1]), .Out(multi23[21][i23]));
      FP16_Multiply stage022(.A(feature4Weight_22), .B(data_array[j23+4][i23+2]), .Out(multi23[22][i23]));
      FP16_Multiply stage023(.A(feature4Weight_23), .B(data_array[j23+4][i23+3]), .Out(multi23[23][i23]));
      FP16_Multiply stage024(.A(feature4Weight_24), .B(data_array[j23+4][i23+4]), .Out(multi23[24][i23]));
      
      ////Sum Stage 1
      FP16_Add stage025(.A(multi23[0][i23]), .B(multi23[1][i23]), .Out(sum23[0][i23]));
      FP16_Add stage026(.A(multi23[2][i23]), .B(multi23[3][i23]), .Out(sum23[1][i23]));
      FP16_Add stage027(.A(multi23[4][i23]), .B(multi23[5][i23]), .Out(sum23[2][i23]));
      FP16_Add stage028(.A(multi23[6][i23]), .B(multi23[7][i23]), .Out(sum23[3][i23]));
      FP16_Add stage029(.A(multi23[8][i23]), .B(multi23[9][i23]), .Out(sum23[4][i23]));
      FP16_Add stage030(.A(multi23[10][i23]), .B(multi23[11][i23]), .Out(sum23[5][i23]));
      FP16_Add stage031(.A(multi23[12][i23]), .B(multi23[13][i23]), .Out(sum23[6][i23]));
      FP16_Add stage032(.A(multi23[14][i23]), .B(multi23[15][i23]), .Out(sum23[7][i23]));
      FP16_Add stage033(.A(multi23[16][i23]), .B(multi23[17][i23]), .Out(sum23[8][i23]));
      FP16_Add stage034(.A(multi23[18][i23]), .B(multi23[19][i23]), .Out(sum23[9][i23]));
      FP16_Add stage035(.A(multi23[20][i23]), .B(multi23[21][i23]), .Out(sum23[10][i23]));
      FP16_Add stage036(.A(multi23[22][i23]), .B(multi23[23][i23]), .Out(sum23[11][i23]));
      
      ////Sum Stage 2
      FP16_Add stage037(.A(sum23[0][i23]), .B(sum23[1][i23]), .Out(sum23[12][i23]));
      FP16_Add stage038(.A(sum23[2][i23]), .B(sum23[3][i23]), .Out(sum23[13][i23]));
      FP16_Add stage039(.A(sum23[4][i23]), .B(sum23[5][i23]), .Out(sum23[14][i23]));
      FP16_Add stage040(.A(sum23[6][i23]), .B(sum23[7][i23]), .Out(sum23[15][i23]));
      FP16_Add stage041(.A(sum23[8][i23]), .B(sum23[9][i23]), .Out(sum23[16][i23]));
      FP16_Add stage042(.A(sum23[10][i23]), .B(sum23[11][i23]), .Out(sum23[17][i23]));
      
      ////Sum Stage 3
      FP16_Add stage043(.A(sum23[12][i23]), .B(sum23[13][i23]), .Out(sum23[18][i23]));
      FP16_Add stage044(.A(sum23[14][i23]), .B(sum23[15][i23]), .Out(sum23[19][i23]));
      FP16_Add stage045(.A(sum23[16][i23]), .B(sum23[17][i23]), .Out(sum23[20][i23]));
      
      ////Sum Stage 4
      FP16_Add stage046(.A(sum23[18][i23]), .B(sum23[19][i23]), .Out(sum23[21][i23]));
      FP16_Add stage047(.A(sum23[20][i23]), .B(multi23[24][i23]), .Out(sum23[22][i23]));
      
      ////Sum Stage 5
      FP16_Add stage048(.A(sum23[21][i23]), .B(sum23[22][i23]), .Out(sum23[23][i23]));
      
      ////Sum Stage 6
      FP16_Add stage049(.A(sum23[23][i23]), .B(feature4Bias), .Out(data_11_array[j23][i23]));
    end
  endgenerate 
  
  localparam integer c0 = 0;
    generate 
        localparam integer d0 = 0;
        for (n0 = 0; n0 < 16; n0 = n0 + 1) 
        begin: outbit0
            assign data_11[n0 + d0*16 + c0*28*16] = data_11_array[c0][d0][n0];
        end
    endgenerate
    generate 
        localparam integer d1 = 1;
        for (n1 = 0; n1 < 16; n1 = n1 + 1) 
        begin: outbit1
            assign data_11[n1 + d1*16 + c0*28*16] = data_11_array[c0][d1][n1];
        end
    endgenerate
    generate 
        localparam integer d2 = 2;
        for (n2 = 0; n2 < 16; n2 = n2 + 1) 
        begin: outbit2
            assign data_11[n2 + d2*16 + c0*28*16] = data_11_array[c0][d2][n2];
        end
    endgenerate
    generate 
        localparam integer d3 = 3;
        for (n3 = 0; n3 < 16; n3 = n3 + 1) 
        begin: outbit3
            assign data_11[n3 + d3*16 + c0*28*16] = data_11_array[c0][d3][n3];
        end
    endgenerate
    generate 
        localparam integer d4 = 4;
        for (n4 = 0; n4 < 16; n4 = n4 + 1) 
        begin: outbit4
            assign data_11[n4 + d4*16 + c0*28*16] = data_11_array[c0][d4][n4];
        end
    endgenerate
    generate 
        localparam integer d5 = 5;
        for (n5 = 0; n5 < 16; n5 = n5 + 1) 
        begin: outbit5
            assign data_11[n5 + d5*16 + c0*28*16] = data_11_array[c0][d5][n5];
        end
    endgenerate
    generate 
        localparam integer d6 = 6;
        for (n6 = 0; n6 < 16; n6 = n6 + 1) 
        begin: outbit6
            assign data_11[n6 + d6*16 + c0*28*16] = data_11_array[c0][d6][n6];
        end
    endgenerate
    generate 
        localparam integer d7 = 7;
        for (n7 = 0; n7 < 16; n7 = n7 + 1) 
        begin: outbit7
            assign data_11[n7 + d7*16 + c0*28*16] = data_11_array[c0][d7][n7];
        end
    endgenerate
    generate 
        localparam integer d8 = 8;
        for (n8 = 0; n8 < 16; n8 = n8 + 1) 
        begin: outbit8
            assign data_11[n8 + d8*16 + c0*28*16] = data_11_array[c0][d8][n8];
        end
    endgenerate
    generate 
        localparam integer d9 = 9;
        for (n9 = 0; n9 < 16; n9 = n9 + 1) 
        begin: outbit9
            assign data_11[n9 + d9*16 + c0*28*16] = data_11_array[c0][d9][n9];
        end
    endgenerate
    generate 
        localparam integer d10 = 10;
        for (n10 = 0; n10 < 16; n10 = n10 + 1) 
        begin: outbit10
            assign data_11[n10 + d10*16 + c0*28*16] = data_11_array[c0][d10][n10];
        end
    endgenerate
    generate 
        localparam integer d11 = 11;
        for (n11 = 0; n11 < 16; n11 = n11 + 1) 
        begin: outbit11
            assign data_11[n11 + d11*16 + c0*28*16] = data_11_array[c0][d11][n11];
        end
    endgenerate
    generate 
        localparam integer d12 = 12;
        for (n12 = 0; n12 < 16; n12 = n12 + 1) 
        begin: outbit12
            assign data_11[n12 + d12*16 + c0*28*16] = data_11_array[c0][d12][n12];
        end
    endgenerate
    generate 
        localparam integer d13 = 13;
        for (n13 = 0; n13 < 16; n13 = n13 + 1) 
        begin: outbit13
            assign data_11[n13 + d13*16 + c0*28*16] = data_11_array[c0][d13][n13];
        end
    endgenerate
    generate 
        localparam integer d14 = 14;
        for (n14 = 0; n14 < 16; n14 = n14 + 1) 
        begin: outbit14
            assign data_11[n14 + d14*16 + c0*28*16] = data_11_array[c0][d14][n14];
        end
    endgenerate
    generate 
        localparam integer d15 = 15;
        for (n15 = 0; n15 < 16; n15 = n15 + 1) 
        begin: outbit15
            assign data_11[n15 + d15*16 + c0*28*16] = data_11_array[c0][d15][n15];
        end
    endgenerate
    generate 
        localparam integer d16 = 16;
        for (n16 = 0; n16 < 16; n16 = n16 + 1) 
        begin: outbit16
            assign data_11[n16 + d16*16 + c0*28*16] = data_11_array[c0][d16][n16];
        end
    endgenerate
    generate 
        localparam integer d17 = 17;
        for (n17 = 0; n17 < 16; n17 = n17 + 1) 
        begin: outbit17
            assign data_11[n17 + d17*16 + c0*28*16] = data_11_array[c0][d17][n17];
        end
    endgenerate
    generate 
        localparam integer d18 = 18;
        for (n18 = 0; n18 < 16; n18 = n18 + 1) 
        begin: outbit18
            assign data_11[n18 + d18*16 + c0*28*16] = data_11_array[c0][d18][n18];
        end
    endgenerate
    generate 
        localparam integer d19 = 19;
        for (n19 = 0; n19 < 16; n19 = n19 + 1) 
        begin: outbit19
            assign data_11[n19 + d19*16 + c0*28*16] = data_11_array[c0][d19][n19];
        end
    endgenerate
    generate 
        localparam integer d20 = 20;
        for (n20 = 0; n20 < 16; n20 = n20 + 1) 
        begin: outbit20
            assign data_11[n20 + d20*16 + c0*28*16] = data_11_array[c0][d20][n20];
        end
    endgenerate
    generate 
        localparam integer d21 = 21;
        for (n21 = 0; n21 < 16; n21 = n21 + 1) 
        begin: outbit21
            assign data_11[n21 + d21*16 + c0*28*16] = data_11_array[c0][d21][n21];
        end
    endgenerate
    generate 
        localparam integer d22 = 22;
        for (n22 = 0; n22 < 16; n22 = n22 + 1) 
        begin: outbit22
            assign data_11[n22 + d22*16 + c0*28*16] = data_11_array[c0][d22][n22];
        end
    endgenerate
    generate 
        localparam integer d23 = 23;
        for (n23 = 0; n23 < 16; n23 = n23 + 1) 
        begin: outbit23
            assign data_11[n23 + d23*16 + c0*28*16] = data_11_array[c0][d23][n23];
        end
    endgenerate
    generate 
        localparam integer d24 = 24;
        for (n24 = 0; n24 < 16; n24 = n24 + 1) 
        begin: outbit24
            assign data_11[n24 + d24*16 + c0*28*16] = data_11_array[c0][d24][n24];
        end
    endgenerate
    generate 
        localparam integer d25 = 25;
        for (n25 = 0; n25 < 16; n25 = n25 + 1) 
        begin: outbit25
            assign data_11[n25 + d25*16 + c0*28*16] = data_11_array[c0][d25][n25];
        end
    endgenerate
    generate 
        localparam integer d26 = 26;
        for (n26 = 0; n26 < 16; n26 = n26 + 1) 
        begin: outbit26
            assign data_11[n26 + d26*16 + c0*28*16] = data_11_array[c0][d26][n26];
        end
    endgenerate
    generate 
        localparam integer d27 = 27;
        for (n27 = 0; n27 < 16; n27 = n27 + 1) 
        begin: outbit27
            assign data_11[n27 + d27*16 + c0*28*16] = data_11_array[c0][d27][n27];
        end
    endgenerate
    localparam integer c1 = 1;
    generate 
        localparam integer d28 = 0;
        for (n28 = 0; n28 < 16; n28 = n28 + 1) 
        begin: outbit28
            assign data_11[n28 + d28*16 + c1*28*16] = data_11_array[c1][d28][n28];
        end
    endgenerate
    generate 
        localparam integer d29 = 1;
        for (n29 = 0; n29 < 16; n29 = n29 + 1) 
        begin: outbit29
            assign data_11[n29 + d29*16 + c1*28*16] = data_11_array[c1][d29][n29];
        end
    endgenerate
    generate 
        localparam integer d30 = 2;
        for (n30 = 0; n30 < 16; n30 = n30 + 1) 
        begin: outbit30
            assign data_11[n30 + d30*16 + c1*28*16] = data_11_array[c1][d30][n30];
        end
    endgenerate
    generate 
        localparam integer d31 = 3;
        for (n31 = 0; n31 < 16; n31 = n31 + 1) 
        begin: outbit31
            assign data_11[n31 + d31*16 + c1*28*16] = data_11_array[c1][d31][n31];
        end
    endgenerate
    generate 
        localparam integer d32 = 4;
        for (n32 = 0; n32 < 16; n32 = n32 + 1) 
        begin: outbit32
            assign data_11[n32 + d32*16 + c1*28*16] = data_11_array[c1][d32][n32];
        end
    endgenerate
    generate 
        localparam integer d33 = 5;
        for (n33 = 0; n33 < 16; n33 = n33 + 1) 
        begin: outbit33
            assign data_11[n33 + d33*16 + c1*28*16] = data_11_array[c1][d33][n33];
        end
    endgenerate
    generate 
        localparam integer d34 = 6;
        for (n34 = 0; n34 < 16; n34 = n34 + 1) 
        begin: outbit34
            assign data_11[n34 + d34*16 + c1*28*16] = data_11_array[c1][d34][n34];
        end
    endgenerate
    generate 
        localparam integer d35 = 7;
        for (n35 = 0; n35 < 16; n35 = n35 + 1) 
        begin: outbit35
            assign data_11[n35 + d35*16 + c1*28*16] = data_11_array[c1][d35][n35];
        end
    endgenerate
    generate 
        localparam integer d36 = 8;
        for (n36 = 0; n36 < 16; n36 = n36 + 1) 
        begin: outbit36
            assign data_11[n36 + d36*16 + c1*28*16] = data_11_array[c1][d36][n36];
        end
    endgenerate
    generate 
        localparam integer d37 = 9;
        for (n37 = 0; n37 < 16; n37 = n37 + 1) 
        begin: outbit37
            assign data_11[n37 + d37*16 + c1*28*16] = data_11_array[c1][d37][n37];
        end
    endgenerate
    generate 
        localparam integer d38 = 10;
        for (n38 = 0; n38 < 16; n38 = n38 + 1) 
        begin: outbit38
            assign data_11[n38 + d38*16 + c1*28*16] = data_11_array[c1][d38][n38];
        end
    endgenerate
    generate 
        localparam integer d39 = 11;
        for (n39 = 0; n39 < 16; n39 = n39 + 1) 
        begin: outbit39
            assign data_11[n39 + d39*16 + c1*28*16] = data_11_array[c1][d39][n39];
        end
    endgenerate
    generate 
        localparam integer d40 = 12;
        for (n40 = 0; n40 < 16; n40 = n40 + 1) 
        begin: outbit40
            assign data_11[n40 + d40*16 + c1*28*16] = data_11_array[c1][d40][n40];
        end
    endgenerate
    generate 
        localparam integer d41 = 13;
        for (n41 = 0; n41 < 16; n41 = n41 + 1) 
        begin: outbit41
            assign data_11[n41 + d41*16 + c1*28*16] = data_11_array[c1][d41][n41];
        end
    endgenerate
    generate 
        localparam integer d42 = 14;
        for (n42 = 0; n42 < 16; n42 = n42 + 1) 
        begin: outbit42
            assign data_11[n42 + d42*16 + c1*28*16] = data_11_array[c1][d42][n42];
        end
    endgenerate
    generate 
        localparam integer d43 = 15;
        for (n43 = 0; n43 < 16; n43 = n43 + 1) 
        begin: outbit43
            assign data_11[n43 + d43*16 + c1*28*16] = data_11_array[c1][d43][n43];
        end
    endgenerate
    generate 
        localparam integer d44 = 16;
        for (n44 = 0; n44 < 16; n44 = n44 + 1) 
        begin: outbit44
            assign data_11[n44 + d44*16 + c1*28*16] = data_11_array[c1][d44][n44];
        end
    endgenerate
    generate 
        localparam integer d45 = 17;
        for (n45 = 0; n45 < 16; n45 = n45 + 1) 
        begin: outbit45
            assign data_11[n45 + d45*16 + c1*28*16] = data_11_array[c1][d45][n45];
        end
    endgenerate
    generate 
        localparam integer d46 = 18;
        for (n46 = 0; n46 < 16; n46 = n46 + 1) 
        begin: outbit46
            assign data_11[n46 + d46*16 + c1*28*16] = data_11_array[c1][d46][n46];
        end
    endgenerate
    generate 
        localparam integer d47 = 19;
        for (n47 = 0; n47 < 16; n47 = n47 + 1) 
        begin: outbit47
            assign data_11[n47 + d47*16 + c1*28*16] = data_11_array[c1][d47][n47];
        end
    endgenerate
    generate 
        localparam integer d48 = 20;
        for (n48 = 0; n48 < 16; n48 = n48 + 1) 
        begin: outbit48
            assign data_11[n48 + d48*16 + c1*28*16] = data_11_array[c1][d48][n48];
        end
    endgenerate
    generate 
        localparam integer d49 = 21;
        for (n49 = 0; n49 < 16; n49 = n49 + 1) 
        begin: outbit49
            assign data_11[n49 + d49*16 + c1*28*16] = data_11_array[c1][d49][n49];
        end
    endgenerate
    generate 
        localparam integer d50 = 22;
        for (n50 = 0; n50 < 16; n50 = n50 + 1) 
        begin: outbit50
            assign data_11[n50 + d50*16 + c1*28*16] = data_11_array[c1][d50][n50];
        end
    endgenerate
    generate 
        localparam integer d51 = 23;
        for (n51 = 0; n51 < 16; n51 = n51 + 1) 
        begin: outbit51
            assign data_11[n51 + d51*16 + c1*28*16] = data_11_array[c1][d51][n51];
        end
    endgenerate
    generate 
        localparam integer d52 = 24;
        for (n52 = 0; n52 < 16; n52 = n52 + 1) 
        begin: outbit52
            assign data_11[n52 + d52*16 + c1*28*16] = data_11_array[c1][d52][n52];
        end
    endgenerate
    generate 
        localparam integer d53 = 25;
        for (n53 = 0; n53 < 16; n53 = n53 + 1) 
        begin: outbit53
            assign data_11[n53 + d53*16 + c1*28*16] = data_11_array[c1][d53][n53];
        end
    endgenerate
    generate 
        localparam integer d54 = 26;
        for (n54 = 0; n54 < 16; n54 = n54 + 1) 
        begin: outbit54
            assign data_11[n54 + d54*16 + c1*28*16] = data_11_array[c1][d54][n54];
        end
    endgenerate
    generate 
        localparam integer d55 = 27;
        for (n55 = 0; n55 < 16; n55 = n55 + 1) 
        begin: outbit55
            assign data_11[n55 + d55*16 + c1*28*16] = data_11_array[c1][d55][n55];
        end
    endgenerate
    localparam integer c2 = 2;
    generate 
        localparam integer d56 = 0;
        for (n56 = 0; n56 < 16; n56 = n56 + 1) 
        begin: outbit56
            assign data_11[n56 + d56*16 + c2*28*16] = data_11_array[c2][d56][n56];
        end
    endgenerate
    generate 
        localparam integer d57 = 1;
        for (n57 = 0; n57 < 16; n57 = n57 + 1) 
        begin: outbit57
            assign data_11[n57 + d57*16 + c2*28*16] = data_11_array[c2][d57][n57];
        end
    endgenerate
    generate 
        localparam integer d58 = 2;
        for (n58 = 0; n58 < 16; n58 = n58 + 1) 
        begin: outbit58
            assign data_11[n58 + d58*16 + c2*28*16] = data_11_array[c2][d58][n58];
        end
    endgenerate
    generate 
        localparam integer d59 = 3;
        for (n59 = 0; n59 < 16; n59 = n59 + 1) 
        begin: outbit59
            assign data_11[n59 + d59*16 + c2*28*16] = data_11_array[c2][d59][n59];
        end
    endgenerate
    generate 
        localparam integer d60 = 4;
        for (n60 = 0; n60 < 16; n60 = n60 + 1) 
        begin: outbit60
            assign data_11[n60 + d60*16 + c2*28*16] = data_11_array[c2][d60][n60];
        end
    endgenerate
    generate 
        localparam integer d61 = 5;
        for (n61 = 0; n61 < 16; n61 = n61 + 1) 
        begin: outbit61
            assign data_11[n61 + d61*16 + c2*28*16] = data_11_array[c2][d61][n61];
        end
    endgenerate
    generate 
        localparam integer d62 = 6;
        for (n62 = 0; n62 < 16; n62 = n62 + 1) 
        begin: outbit62
            assign data_11[n62 + d62*16 + c2*28*16] = data_11_array[c2][d62][n62];
        end
    endgenerate
    generate 
        localparam integer d63 = 7;
        for (n63 = 0; n63 < 16; n63 = n63 + 1) 
        begin: outbit63
            assign data_11[n63 + d63*16 + c2*28*16] = data_11_array[c2][d63][n63];
        end
    endgenerate
    generate 
        localparam integer d64 = 8;
        for (n64 = 0; n64 < 16; n64 = n64 + 1) 
        begin: outbit64
            assign data_11[n64 + d64*16 + c2*28*16] = data_11_array[c2][d64][n64];
        end
    endgenerate
    generate 
        localparam integer d65 = 9;
        for (n65 = 0; n65 < 16; n65 = n65 + 1) 
        begin: outbit65
            assign data_11[n65 + d65*16 + c2*28*16] = data_11_array[c2][d65][n65];
        end
    endgenerate
    generate 
        localparam integer d66 = 10;
        for (n66 = 0; n66 < 16; n66 = n66 + 1) 
        begin: outbit66
            assign data_11[n66 + d66*16 + c2*28*16] = data_11_array[c2][d66][n66];
        end
    endgenerate
    generate 
        localparam integer d67 = 11;
        for (n67 = 0; n67 < 16; n67 = n67 + 1) 
        begin: outbit67
            assign data_11[n67 + d67*16 + c2*28*16] = data_11_array[c2][d67][n67];
        end
    endgenerate
    generate 
        localparam integer d68 = 12;
        for (n68 = 0; n68 < 16; n68 = n68 + 1) 
        begin: outbit68
            assign data_11[n68 + d68*16 + c2*28*16] = data_11_array[c2][d68][n68];
        end
    endgenerate
    generate 
        localparam integer d69 = 13;
        for (n69 = 0; n69 < 16; n69 = n69 + 1) 
        begin: outbit69
            assign data_11[n69 + d69*16 + c2*28*16] = data_11_array[c2][d69][n69];
        end
    endgenerate
    generate 
        localparam integer d70 = 14;
        for (n70 = 0; n70 < 16; n70 = n70 + 1) 
        begin: outbit70
            assign data_11[n70 + d70*16 + c2*28*16] = data_11_array[c2][d70][n70];
        end
    endgenerate
    generate 
        localparam integer d71 = 15;
        for (n71 = 0; n71 < 16; n71 = n71 + 1) 
        begin: outbit71
            assign data_11[n71 + d71*16 + c2*28*16] = data_11_array[c2][d71][n71];
        end
    endgenerate
    generate 
        localparam integer d72 = 16;
        for (n72 = 0; n72 < 16; n72 = n72 + 1) 
        begin: outbit72
            assign data_11[n72 + d72*16 + c2*28*16] = data_11_array[c2][d72][n72];
        end
    endgenerate
    generate 
        localparam integer d73 = 17;
        for (n73 = 0; n73 < 16; n73 = n73 + 1) 
        begin: outbit73
            assign data_11[n73 + d73*16 + c2*28*16] = data_11_array[c2][d73][n73];
        end
    endgenerate
    generate 
        localparam integer d74 = 18;
        for (n74 = 0; n74 < 16; n74 = n74 + 1) 
        begin: outbit74
            assign data_11[n74 + d74*16 + c2*28*16] = data_11_array[c2][d74][n74];
        end
    endgenerate
    generate 
        localparam integer d75 = 19;
        for (n75 = 0; n75 < 16; n75 = n75 + 1) 
        begin: outbit75
            assign data_11[n75 + d75*16 + c2*28*16] = data_11_array[c2][d75][n75];
        end
    endgenerate
    generate 
        localparam integer d76 = 20;
        for (n76 = 0; n76 < 16; n76 = n76 + 1) 
        begin: outbit76
            assign data_11[n76 + d76*16 + c2*28*16] = data_11_array[c2][d76][n76];
        end
    endgenerate
    generate 
        localparam integer d77 = 21;
        for (n77 = 0; n77 < 16; n77 = n77 + 1) 
        begin: outbit77
            assign data_11[n77 + d77*16 + c2*28*16] = data_11_array[c2][d77][n77];
        end
    endgenerate
    generate 
        localparam integer d78 = 22;
        for (n78 = 0; n78 < 16; n78 = n78 + 1) 
        begin: outbit78
            assign data_11[n78 + d78*16 + c2*28*16] = data_11_array[c2][d78][n78];
        end
    endgenerate
    generate 
        localparam integer d79 = 23;
        for (n79 = 0; n79 < 16; n79 = n79 + 1) 
        begin: outbit79
            assign data_11[n79 + d79*16 + c2*28*16] = data_11_array[c2][d79][n79];
        end
    endgenerate
    generate 
        localparam integer d80 = 24;
        for (n80 = 0; n80 < 16; n80 = n80 + 1) 
        begin: outbit80
            assign data_11[n80 + d80*16 + c2*28*16] = data_11_array[c2][d80][n80];
        end
    endgenerate
    generate 
        localparam integer d81 = 25;
        for (n81 = 0; n81 < 16; n81 = n81 + 1) 
        begin: outbit81
            assign data_11[n81 + d81*16 + c2*28*16] = data_11_array[c2][d81][n81];
        end
    endgenerate
    generate 
        localparam integer d82 = 26;
        for (n82 = 0; n82 < 16; n82 = n82 + 1) 
        begin: outbit82
            assign data_11[n82 + d82*16 + c2*28*16] = data_11_array[c2][d82][n82];
        end
    endgenerate
    generate 
        localparam integer d83 = 27;
        for (n83 = 0; n83 < 16; n83 = n83 + 1) 
        begin: outbit83
            assign data_11[n83 + d83*16 + c2*28*16] = data_11_array[c2][d83][n83];
        end
    endgenerate
    localparam integer c3 = 3;
    generate 
        localparam integer d84 = 0;
        for (n84 = 0; n84 < 16; n84 = n84 + 1) 
        begin: outbit84
            assign data_11[n84 + d84*16 + c3*28*16] = data_11_array[c3][d84][n84];
        end
    endgenerate
    generate 
        localparam integer d85 = 1;
        for (n85 = 0; n85 < 16; n85 = n85 + 1) 
        begin: outbit85
            assign data_11[n85 + d85*16 + c3*28*16] = data_11_array[c3][d85][n85];
        end
    endgenerate
    generate 
        localparam integer d86 = 2;
        for (n86 = 0; n86 < 16; n86 = n86 + 1) 
        begin: outbit86
            assign data_11[n86 + d86*16 + c3*28*16] = data_11_array[c3][d86][n86];
        end
    endgenerate
    generate 
        localparam integer d87 = 3;
        for (n87 = 0; n87 < 16; n87 = n87 + 1) 
        begin: outbit87
            assign data_11[n87 + d87*16 + c3*28*16] = data_11_array[c3][d87][n87];
        end
    endgenerate
    generate 
        localparam integer d88 = 4;
        for (n88 = 0; n88 < 16; n88 = n88 + 1) 
        begin: outbit88
            assign data_11[n88 + d88*16 + c3*28*16] = data_11_array[c3][d88][n88];
        end
    endgenerate
    generate 
        localparam integer d89 = 5;
        for (n89 = 0; n89 < 16; n89 = n89 + 1) 
        begin: outbit89
            assign data_11[n89 + d89*16 + c3*28*16] = data_11_array[c3][d89][n89];
        end
    endgenerate
    generate 
        localparam integer d90 = 6;
        for (n90 = 0; n90 < 16; n90 = n90 + 1) 
        begin: outbit90
            assign data_11[n90 + d90*16 + c3*28*16] = data_11_array[c3][d90][n90];
        end
    endgenerate
    generate 
        localparam integer d91 = 7;
        for (n91 = 0; n91 < 16; n91 = n91 + 1) 
        begin: outbit91
            assign data_11[n91 + d91*16 + c3*28*16] = data_11_array[c3][d91][n91];
        end
    endgenerate
    generate 
        localparam integer d92 = 8;
        for (n92 = 0; n92 < 16; n92 = n92 + 1) 
        begin: outbit92
            assign data_11[n92 + d92*16 + c3*28*16] = data_11_array[c3][d92][n92];
        end
    endgenerate
    generate 
        localparam integer d93 = 9;
        for (n93 = 0; n93 < 16; n93 = n93 + 1) 
        begin: outbit93
            assign data_11[n93 + d93*16 + c3*28*16] = data_11_array[c3][d93][n93];
        end
    endgenerate
    generate 
        localparam integer d94 = 10;
        for (n94 = 0; n94 < 16; n94 = n94 + 1) 
        begin: outbit94
            assign data_11[n94 + d94*16 + c3*28*16] = data_11_array[c3][d94][n94];
        end
    endgenerate
    generate 
        localparam integer d95 = 11;
        for (n95 = 0; n95 < 16; n95 = n95 + 1) 
        begin: outbit95
            assign data_11[n95 + d95*16 + c3*28*16] = data_11_array[c3][d95][n95];
        end
    endgenerate
    generate 
        localparam integer d96 = 12;
        for (n96 = 0; n96 < 16; n96 = n96 + 1) 
        begin: outbit96
            assign data_11[n96 + d96*16 + c3*28*16] = data_11_array[c3][d96][n96];
        end
    endgenerate
    generate 
        localparam integer d97 = 13;
        for (n97 = 0; n97 < 16; n97 = n97 + 1) 
        begin: outbit97
            assign data_11[n97 + d97*16 + c3*28*16] = data_11_array[c3][d97][n97];
        end
    endgenerate
    generate 
        localparam integer d98 = 14;
        for (n98 = 0; n98 < 16; n98 = n98 + 1) 
        begin: outbit98
            assign data_11[n98 + d98*16 + c3*28*16] = data_11_array[c3][d98][n98];
        end
    endgenerate
    generate 
        localparam integer d99 = 15;
        for (n99 = 0; n99 < 16; n99 = n99 + 1) 
        begin: outbit99
            assign data_11[n99 + d99*16 + c3*28*16] = data_11_array[c3][d99][n99];
        end
    endgenerate
    generate 
        localparam integer d100 = 16;
        for (n100 = 0; n100 < 16; n100 = n100 + 1) 
        begin: outbit100
            assign data_11[n100 + d100*16 + c3*28*16] = data_11_array[c3][d100][n100];
        end
    endgenerate
    generate 
        localparam integer d101 = 17;
        for (n101 = 0; n101 < 16; n101 = n101 + 1) 
        begin: outbit101
            assign data_11[n101 + d101*16 + c3*28*16] = data_11_array[c3][d101][n101];
        end
    endgenerate
    generate 
        localparam integer d102 = 18;
        for (n102 = 0; n102 < 16; n102 = n102 + 1) 
        begin: outbit102
            assign data_11[n102 + d102*16 + c3*28*16] = data_11_array[c3][d102][n102];
        end
    endgenerate
    generate 
        localparam integer d103 = 19;
        for (n103 = 0; n103 < 16; n103 = n103 + 1) 
        begin: outbit103
            assign data_11[n103 + d103*16 + c3*28*16] = data_11_array[c3][d103][n103];
        end
    endgenerate
    generate 
        localparam integer d104 = 20;
        for (n104 = 0; n104 < 16; n104 = n104 + 1) 
        begin: outbit104
            assign data_11[n104 + d104*16 + c3*28*16] = data_11_array[c3][d104][n104];
        end
    endgenerate
    generate 
        localparam integer d105 = 21;
        for (n105 = 0; n105 < 16; n105 = n105 + 1) 
        begin: outbit105
            assign data_11[n105 + d105*16 + c3*28*16] = data_11_array[c3][d105][n105];
        end
    endgenerate
    generate 
        localparam integer d106 = 22;
        for (n106 = 0; n106 < 16; n106 = n106 + 1) 
        begin: outbit106
            assign data_11[n106 + d106*16 + c3*28*16] = data_11_array[c3][d106][n106];
        end
    endgenerate
    generate 
        localparam integer d107 = 23;
        for (n107 = 0; n107 < 16; n107 = n107 + 1) 
        begin: outbit107
            assign data_11[n107 + d107*16 + c3*28*16] = data_11_array[c3][d107][n107];
        end
    endgenerate
    generate 
        localparam integer d108 = 24;
        for (n108 = 0; n108 < 16; n108 = n108 + 1) 
        begin: outbit108
            assign data_11[n108 + d108*16 + c3*28*16] = data_11_array[c3][d108][n108];
        end
    endgenerate
    generate 
        localparam integer d109 = 25;
        for (n109 = 0; n109 < 16; n109 = n109 + 1) 
        begin: outbit109
            assign data_11[n109 + d109*16 + c3*28*16] = data_11_array[c3][d109][n109];
        end
    endgenerate
    generate 
        localparam integer d110 = 26;
        for (n110 = 0; n110 < 16; n110 = n110 + 1) 
        begin: outbit110
            assign data_11[n110 + d110*16 + c3*28*16] = data_11_array[c3][d110][n110];
        end
    endgenerate
    generate 
        localparam integer d111 = 27;
        for (n111 = 0; n111 < 16; n111 = n111 + 1) 
        begin: outbit111
            assign data_11[n111 + d111*16 + c3*28*16] = data_11_array[c3][d111][n111];
        end
    endgenerate
    localparam integer c4 = 4;
    generate 
        localparam integer d112 = 0;
        for (n112 = 0; n112 < 16; n112 = n112 + 1) 
        begin: outbit112
            assign data_11[n112 + d112*16 + c4*28*16] = data_11_array[c4][d112][n112];
        end
    endgenerate
    generate 
        localparam integer d113 = 1;
        for (n113 = 0; n113 < 16; n113 = n113 + 1) 
        begin: outbit113
            assign data_11[n113 + d113*16 + c4*28*16] = data_11_array[c4][d113][n113];
        end
    endgenerate
    generate 
        localparam integer d114 = 2;
        for (n114 = 0; n114 < 16; n114 = n114 + 1) 
        begin: outbit114
            assign data_11[n114 + d114*16 + c4*28*16] = data_11_array[c4][d114][n114];
        end
    endgenerate
    generate 
        localparam integer d115 = 3;
        for (n115 = 0; n115 < 16; n115 = n115 + 1) 
        begin: outbit115
            assign data_11[n115 + d115*16 + c4*28*16] = data_11_array[c4][d115][n115];
        end
    endgenerate
    generate 
        localparam integer d116 = 4;
        for (n116 = 0; n116 < 16; n116 = n116 + 1) 
        begin: outbit116
            assign data_11[n116 + d116*16 + c4*28*16] = data_11_array[c4][d116][n116];
        end
    endgenerate
    generate 
        localparam integer d117 = 5;
        for (n117 = 0; n117 < 16; n117 = n117 + 1) 
        begin: outbit117
            assign data_11[n117 + d117*16 + c4*28*16] = data_11_array[c4][d117][n117];
        end
    endgenerate
    generate 
        localparam integer d118 = 6;
        for (n118 = 0; n118 < 16; n118 = n118 + 1) 
        begin: outbit118
            assign data_11[n118 + d118*16 + c4*28*16] = data_11_array[c4][d118][n118];
        end
    endgenerate
    generate 
        localparam integer d119 = 7;
        for (n119 = 0; n119 < 16; n119 = n119 + 1) 
        begin: outbit119
            assign data_11[n119 + d119*16 + c4*28*16] = data_11_array[c4][d119][n119];
        end
    endgenerate
    generate 
        localparam integer d120 = 8;
        for (n120 = 0; n120 < 16; n120 = n120 + 1) 
        begin: outbit120
            assign data_11[n120 + d120*16 + c4*28*16] = data_11_array[c4][d120][n120];
        end
    endgenerate
    generate 
        localparam integer d121 = 9;
        for (n121 = 0; n121 < 16; n121 = n121 + 1) 
        begin: outbit121
            assign data_11[n121 + d121*16 + c4*28*16] = data_11_array[c4][d121][n121];
        end
    endgenerate
    generate 
        localparam integer d122 = 10;
        for (n122 = 0; n122 < 16; n122 = n122 + 1) 
        begin: outbit122
            assign data_11[n122 + d122*16 + c4*28*16] = data_11_array[c4][d122][n122];
        end
    endgenerate
    generate 
        localparam integer d123 = 11;
        for (n123 = 0; n123 < 16; n123 = n123 + 1) 
        begin: outbit123
            assign data_11[n123 + d123*16 + c4*28*16] = data_11_array[c4][d123][n123];
        end
    endgenerate
    generate 
        localparam integer d124 = 12;
        for (n124 = 0; n124 < 16; n124 = n124 + 1) 
        begin: outbit124
            assign data_11[n124 + d124*16 + c4*28*16] = data_11_array[c4][d124][n124];
        end
    endgenerate
    generate 
        localparam integer d125 = 13;
        for (n125 = 0; n125 < 16; n125 = n125 + 1) 
        begin: outbit125
            assign data_11[n125 + d125*16 + c4*28*16] = data_11_array[c4][d125][n125];
        end
    endgenerate
    generate 
        localparam integer d126 = 14;
        for (n126 = 0; n126 < 16; n126 = n126 + 1) 
        begin: outbit126
            assign data_11[n126 + d126*16 + c4*28*16] = data_11_array[c4][d126][n126];
        end
    endgenerate
    generate 
        localparam integer d127 = 15;
        for (n127 = 0; n127 < 16; n127 = n127 + 1) 
        begin: outbit127
            assign data_11[n127 + d127*16 + c4*28*16] = data_11_array[c4][d127][n127];
        end
    endgenerate
    generate 
        localparam integer d128 = 16;
        for (n128 = 0; n128 < 16; n128 = n128 + 1) 
        begin: outbit128
            assign data_11[n128 + d128*16 + c4*28*16] = data_11_array[c4][d128][n128];
        end
    endgenerate
    generate 
        localparam integer d129 = 17;
        for (n129 = 0; n129 < 16; n129 = n129 + 1) 
        begin: outbit129
            assign data_11[n129 + d129*16 + c4*28*16] = data_11_array[c4][d129][n129];
        end
    endgenerate
    generate 
        localparam integer d130 = 18;
        for (n130 = 0; n130 < 16; n130 = n130 + 1) 
        begin: outbit130
            assign data_11[n130 + d130*16 + c4*28*16] = data_11_array[c4][d130][n130];
        end
    endgenerate
    generate 
        localparam integer d131 = 19;
        for (n131 = 0; n131 < 16; n131 = n131 + 1) 
        begin: outbit131
            assign data_11[n131 + d131*16 + c4*28*16] = data_11_array[c4][d131][n131];
        end
    endgenerate
    generate 
        localparam integer d132 = 20;
        for (n132 = 0; n132 < 16; n132 = n132 + 1) 
        begin: outbit132
            assign data_11[n132 + d132*16 + c4*28*16] = data_11_array[c4][d132][n132];
        end
    endgenerate
    generate 
        localparam integer d133 = 21;
        for (n133 = 0; n133 < 16; n133 = n133 + 1) 
        begin: outbit133
            assign data_11[n133 + d133*16 + c4*28*16] = data_11_array[c4][d133][n133];
        end
    endgenerate
    generate 
        localparam integer d134 = 22;
        for (n134 = 0; n134 < 16; n134 = n134 + 1) 
        begin: outbit134
            assign data_11[n134 + d134*16 + c4*28*16] = data_11_array[c4][d134][n134];
        end
    endgenerate
    generate 
        localparam integer d135 = 23;
        for (n135 = 0; n135 < 16; n135 = n135 + 1) 
        begin: outbit135
            assign data_11[n135 + d135*16 + c4*28*16] = data_11_array[c4][d135][n135];
        end
    endgenerate
    generate 
        localparam integer d136 = 24;
        for (n136 = 0; n136 < 16; n136 = n136 + 1) 
        begin: outbit136
            assign data_11[n136 + d136*16 + c4*28*16] = data_11_array[c4][d136][n136];
        end
    endgenerate
    generate 
        localparam integer d137 = 25;
        for (n137 = 0; n137 < 16; n137 = n137 + 1) 
        begin: outbit137
            assign data_11[n137 + d137*16 + c4*28*16] = data_11_array[c4][d137][n137];
        end
    endgenerate
    generate 
        localparam integer d138 = 26;
        for (n138 = 0; n138 < 16; n138 = n138 + 1) 
        begin: outbit138
            assign data_11[n138 + d138*16 + c4*28*16] = data_11_array[c4][d138][n138];
        end
    endgenerate
    generate 
        localparam integer d139 = 27;
        for (n139 = 0; n139 < 16; n139 = n139 + 1) 
        begin: outbit139
            assign data_11[n139 + d139*16 + c4*28*16] = data_11_array[c4][d139][n139];
        end
    endgenerate
    localparam integer c5 = 5;
    generate 
        localparam integer d140 = 0;
        for (n140 = 0; n140 < 16; n140 = n140 + 1) 
        begin: outbit140
            assign data_11[n140 + d140*16 + c5*28*16] = data_11_array[c5][d140][n140];
        end
    endgenerate
    generate 
        localparam integer d141 = 1;
        for (n141 = 0; n141 < 16; n141 = n141 + 1) 
        begin: outbit141
            assign data_11[n141 + d141*16 + c5*28*16] = data_11_array[c5][d141][n141];
        end
    endgenerate
    generate 
        localparam integer d142 = 2;
        for (n142 = 0; n142 < 16; n142 = n142 + 1) 
        begin: outbit142
            assign data_11[n142 + d142*16 + c5*28*16] = data_11_array[c5][d142][n142];
        end
    endgenerate
    generate 
        localparam integer d143 = 3;
        for (n143 = 0; n143 < 16; n143 = n143 + 1) 
        begin: outbit143
            assign data_11[n143 + d143*16 + c5*28*16] = data_11_array[c5][d143][n143];
        end
    endgenerate
    generate 
        localparam integer d144 = 4;
        for (n144 = 0; n144 < 16; n144 = n144 + 1) 
        begin: outbit144
            assign data_11[n144 + d144*16 + c5*28*16] = data_11_array[c5][d144][n144];
        end
    endgenerate
    generate 
        localparam integer d145 = 5;
        for (n145 = 0; n145 < 16; n145 = n145 + 1) 
        begin: outbit145
            assign data_11[n145 + d145*16 + c5*28*16] = data_11_array[c5][d145][n145];
        end
    endgenerate
    generate 
        localparam integer d146 = 6;
        for (n146 = 0; n146 < 16; n146 = n146 + 1) 
        begin: outbit146
            assign data_11[n146 + d146*16 + c5*28*16] = data_11_array[c5][d146][n146];
        end
    endgenerate
    generate 
        localparam integer d147 = 7;
        for (n147 = 0; n147 < 16; n147 = n147 + 1) 
        begin: outbit147
            assign data_11[n147 + d147*16 + c5*28*16] = data_11_array[c5][d147][n147];
        end
    endgenerate
    generate 
        localparam integer d148 = 8;
        for (n148 = 0; n148 < 16; n148 = n148 + 1) 
        begin: outbit148
            assign data_11[n148 + d148*16 + c5*28*16] = data_11_array[c5][d148][n148];
        end
    endgenerate
    generate 
        localparam integer d149 = 9;
        for (n149 = 0; n149 < 16; n149 = n149 + 1) 
        begin: outbit149
            assign data_11[n149 + d149*16 + c5*28*16] = data_11_array[c5][d149][n149];
        end
    endgenerate
    generate 
        localparam integer d150 = 10;
        for (n150 = 0; n150 < 16; n150 = n150 + 1) 
        begin: outbit150
            assign data_11[n150 + d150*16 + c5*28*16] = data_11_array[c5][d150][n150];
        end
    endgenerate
    generate 
        localparam integer d151 = 11;
        for (n151 = 0; n151 < 16; n151 = n151 + 1) 
        begin: outbit151
            assign data_11[n151 + d151*16 + c5*28*16] = data_11_array[c5][d151][n151];
        end
    endgenerate
    generate 
        localparam integer d152 = 12;
        for (n152 = 0; n152 < 16; n152 = n152 + 1) 
        begin: outbit152
            assign data_11[n152 + d152*16 + c5*28*16] = data_11_array[c5][d152][n152];
        end
    endgenerate
    generate 
        localparam integer d153 = 13;
        for (n153 = 0; n153 < 16; n153 = n153 + 1) 
        begin: outbit153
            assign data_11[n153 + d153*16 + c5*28*16] = data_11_array[c5][d153][n153];
        end
    endgenerate
    generate 
        localparam integer d154 = 14;
        for (n154 = 0; n154 < 16; n154 = n154 + 1) 
        begin: outbit154
            assign data_11[n154 + d154*16 + c5*28*16] = data_11_array[c5][d154][n154];
        end
    endgenerate
    generate 
        localparam integer d155 = 15;
        for (n155 = 0; n155 < 16; n155 = n155 + 1) 
        begin: outbit155
            assign data_11[n155 + d155*16 + c5*28*16] = data_11_array[c5][d155][n155];
        end
    endgenerate
    generate 
        localparam integer d156 = 16;
        for (n156 = 0; n156 < 16; n156 = n156 + 1) 
        begin: outbit156
            assign data_11[n156 + d156*16 + c5*28*16] = data_11_array[c5][d156][n156];
        end
    endgenerate
    generate 
        localparam integer d157 = 17;
        for (n157 = 0; n157 < 16; n157 = n157 + 1) 
        begin: outbit157
            assign data_11[n157 + d157*16 + c5*28*16] = data_11_array[c5][d157][n157];
        end
    endgenerate
    generate 
        localparam integer d158 = 18;
        for (n158 = 0; n158 < 16; n158 = n158 + 1) 
        begin: outbit158
            assign data_11[n158 + d158*16 + c5*28*16] = data_11_array[c5][d158][n158];
        end
    endgenerate
    generate 
        localparam integer d159 = 19;
        for (n159 = 0; n159 < 16; n159 = n159 + 1) 
        begin: outbit159
            assign data_11[n159 + d159*16 + c5*28*16] = data_11_array[c5][d159][n159];
        end
    endgenerate
    generate 
        localparam integer d160 = 20;
        for (n160 = 0; n160 < 16; n160 = n160 + 1) 
        begin: outbit160
            assign data_11[n160 + d160*16 + c5*28*16] = data_11_array[c5][d160][n160];
        end
    endgenerate
    generate 
        localparam integer d161 = 21;
        for (n161 = 0; n161 < 16; n161 = n161 + 1) 
        begin: outbit161
            assign data_11[n161 + d161*16 + c5*28*16] = data_11_array[c5][d161][n161];
        end
    endgenerate
    generate 
        localparam integer d162 = 22;
        for (n162 = 0; n162 < 16; n162 = n162 + 1) 
        begin: outbit162
            assign data_11[n162 + d162*16 + c5*28*16] = data_11_array[c5][d162][n162];
        end
    endgenerate
    generate 
        localparam integer d163 = 23;
        for (n163 = 0; n163 < 16; n163 = n163 + 1) 
        begin: outbit163
            assign data_11[n163 + d163*16 + c5*28*16] = data_11_array[c5][d163][n163];
        end
    endgenerate
    generate 
        localparam integer d164 = 24;
        for (n164 = 0; n164 < 16; n164 = n164 + 1) 
        begin: outbit164
            assign data_11[n164 + d164*16 + c5*28*16] = data_11_array[c5][d164][n164];
        end
    endgenerate
    generate 
        localparam integer d165 = 25;
        for (n165 = 0; n165 < 16; n165 = n165 + 1) 
        begin: outbit165
            assign data_11[n165 + d165*16 + c5*28*16] = data_11_array[c5][d165][n165];
        end
    endgenerate
    generate 
        localparam integer d166 = 26;
        for (n166 = 0; n166 < 16; n166 = n166 + 1) 
        begin: outbit166
            assign data_11[n166 + d166*16 + c5*28*16] = data_11_array[c5][d166][n166];
        end
    endgenerate
    generate 
        localparam integer d167 = 27;
        for (n167 = 0; n167 < 16; n167 = n167 + 1) 
        begin: outbit167
            assign data_11[n167 + d167*16 + c5*28*16] = data_11_array[c5][d167][n167];
        end
    endgenerate
    localparam integer c6 = 6;
    generate 
        localparam integer d168 = 0;
        for (n168 = 0; n168 < 16; n168 = n168 + 1) 
        begin: outbit168
            assign data_11[n168 + d168*16 + c6*28*16] = data_11_array[c6][d168][n168];
        end
    endgenerate
    generate 
        localparam integer d169 = 1;
        for (n169 = 0; n169 < 16; n169 = n169 + 1) 
        begin: outbit169
            assign data_11[n169 + d169*16 + c6*28*16] = data_11_array[c6][d169][n169];
        end
    endgenerate
    generate 
        localparam integer d170 = 2;
        for (n170 = 0; n170 < 16; n170 = n170 + 1) 
        begin: outbit170
            assign data_11[n170 + d170*16 + c6*28*16] = data_11_array[c6][d170][n170];
        end
    endgenerate
    generate 
        localparam integer d171 = 3;
        for (n171 = 0; n171 < 16; n171 = n171 + 1) 
        begin: outbit171
            assign data_11[n171 + d171*16 + c6*28*16] = data_11_array[c6][d171][n171];
        end
    endgenerate
    generate 
        localparam integer d172 = 4;
        for (n172 = 0; n172 < 16; n172 = n172 + 1) 
        begin: outbit172
            assign data_11[n172 + d172*16 + c6*28*16] = data_11_array[c6][d172][n172];
        end
    endgenerate
    generate 
        localparam integer d173 = 5;
        for (n173 = 0; n173 < 16; n173 = n173 + 1) 
        begin: outbit173
            assign data_11[n173 + d173*16 + c6*28*16] = data_11_array[c6][d173][n173];
        end
    endgenerate
    generate 
        localparam integer d174 = 6;
        for (n174 = 0; n174 < 16; n174 = n174 + 1) 
        begin: outbit174
            assign data_11[n174 + d174*16 + c6*28*16] = data_11_array[c6][d174][n174];
        end
    endgenerate
    generate 
        localparam integer d175 = 7;
        for (n175 = 0; n175 < 16; n175 = n175 + 1) 
        begin: outbit175
            assign data_11[n175 + d175*16 + c6*28*16] = data_11_array[c6][d175][n175];
        end
    endgenerate
    generate 
        localparam integer d176 = 8;
        for (n176 = 0; n176 < 16; n176 = n176 + 1) 
        begin: outbit176
            assign data_11[n176 + d176*16 + c6*28*16] = data_11_array[c6][d176][n176];
        end
    endgenerate
    generate 
        localparam integer d177 = 9;
        for (n177 = 0; n177 < 16; n177 = n177 + 1) 
        begin: outbit177
            assign data_11[n177 + d177*16 + c6*28*16] = data_11_array[c6][d177][n177];
        end
    endgenerate
    generate 
        localparam integer d178 = 10;
        for (n178 = 0; n178 < 16; n178 = n178 + 1) 
        begin: outbit178
            assign data_11[n178 + d178*16 + c6*28*16] = data_11_array[c6][d178][n178];
        end
    endgenerate
    generate 
        localparam integer d179 = 11;
        for (n179 = 0; n179 < 16; n179 = n179 + 1) 
        begin: outbit179
            assign data_11[n179 + d179*16 + c6*28*16] = data_11_array[c6][d179][n179];
        end
    endgenerate
    generate 
        localparam integer d180 = 12;
        for (n180 = 0; n180 < 16; n180 = n180 + 1) 
        begin: outbit180
            assign data_11[n180 + d180*16 + c6*28*16] = data_11_array[c6][d180][n180];
        end
    endgenerate
    generate 
        localparam integer d181 = 13;
        for (n181 = 0; n181 < 16; n181 = n181 + 1) 
        begin: outbit181
            assign data_11[n181 + d181*16 + c6*28*16] = data_11_array[c6][d181][n181];
        end
    endgenerate
    generate 
        localparam integer d182 = 14;
        for (n182 = 0; n182 < 16; n182 = n182 + 1) 
        begin: outbit182
            assign data_11[n182 + d182*16 + c6*28*16] = data_11_array[c6][d182][n182];
        end
    endgenerate
    generate 
        localparam integer d183 = 15;
        for (n183 = 0; n183 < 16; n183 = n183 + 1) 
        begin: outbit183
            assign data_11[n183 + d183*16 + c6*28*16] = data_11_array[c6][d183][n183];
        end
    endgenerate
    generate 
        localparam integer d184 = 16;
        for (n184 = 0; n184 < 16; n184 = n184 + 1) 
        begin: outbit184
            assign data_11[n184 + d184*16 + c6*28*16] = data_11_array[c6][d184][n184];
        end
    endgenerate
    generate 
        localparam integer d185 = 17;
        for (n185 = 0; n185 < 16; n185 = n185 + 1) 
        begin: outbit185
            assign data_11[n185 + d185*16 + c6*28*16] = data_11_array[c6][d185][n185];
        end
    endgenerate
    generate 
        localparam integer d186 = 18;
        for (n186 = 0; n186 < 16; n186 = n186 + 1) 
        begin: outbit186
            assign data_11[n186 + d186*16 + c6*28*16] = data_11_array[c6][d186][n186];
        end
    endgenerate
    generate 
        localparam integer d187 = 19;
        for (n187 = 0; n187 < 16; n187 = n187 + 1) 
        begin: outbit187
            assign data_11[n187 + d187*16 + c6*28*16] = data_11_array[c6][d187][n187];
        end
    endgenerate
    generate 
        localparam integer d188 = 20;
        for (n188 = 0; n188 < 16; n188 = n188 + 1) 
        begin: outbit188
            assign data_11[n188 + d188*16 + c6*28*16] = data_11_array[c6][d188][n188];
        end
    endgenerate
    generate 
        localparam integer d189 = 21;
        for (n189 = 0; n189 < 16; n189 = n189 + 1) 
        begin: outbit189
            assign data_11[n189 + d189*16 + c6*28*16] = data_11_array[c6][d189][n189];
        end
    endgenerate
    generate 
        localparam integer d190 = 22;
        for (n190 = 0; n190 < 16; n190 = n190 + 1) 
        begin: outbit190
            assign data_11[n190 + d190*16 + c6*28*16] = data_11_array[c6][d190][n190];
        end
    endgenerate
    generate 
        localparam integer d191 = 23;
        for (n191 = 0; n191 < 16; n191 = n191 + 1) 
        begin: outbit191
            assign data_11[n191 + d191*16 + c6*28*16] = data_11_array[c6][d191][n191];
        end
    endgenerate
    generate 
        localparam integer d192 = 24;
        for (n192 = 0; n192 < 16; n192 = n192 + 1) 
        begin: outbit192
            assign data_11[n192 + d192*16 + c6*28*16] = data_11_array[c6][d192][n192];
        end
    endgenerate
    generate 
        localparam integer d193 = 25;
        for (n193 = 0; n193 < 16; n193 = n193 + 1) 
        begin: outbit193
            assign data_11[n193 + d193*16 + c6*28*16] = data_11_array[c6][d193][n193];
        end
    endgenerate
    generate 
        localparam integer d194 = 26;
        for (n194 = 0; n194 < 16; n194 = n194 + 1) 
        begin: outbit194
            assign data_11[n194 + d194*16 + c6*28*16] = data_11_array[c6][d194][n194];
        end
    endgenerate
    generate 
        localparam integer d195 = 27;
        for (n195 = 0; n195 < 16; n195 = n195 + 1) 
        begin: outbit195
            assign data_11[n195 + d195*16 + c6*28*16] = data_11_array[c6][d195][n195];
        end
    endgenerate
    localparam integer c7 = 7;
    generate 
        localparam integer d196 = 0;
        for (n196 = 0; n196 < 16; n196 = n196 + 1) 
        begin: outbit196
            assign data_11[n196 + d196*16 + c7*28*16] = data_11_array[c7][d196][n196];
        end
    endgenerate
    generate 
        localparam integer d197 = 1;
        for (n197 = 0; n197 < 16; n197 = n197 + 1) 
        begin: outbit197
            assign data_11[n197 + d197*16 + c7*28*16] = data_11_array[c7][d197][n197];
        end
    endgenerate
    generate 
        localparam integer d198 = 2;
        for (n198 = 0; n198 < 16; n198 = n198 + 1) 
        begin: outbit198
            assign data_11[n198 + d198*16 + c7*28*16] = data_11_array[c7][d198][n198];
        end
    endgenerate
    generate 
        localparam integer d199 = 3;
        for (n199 = 0; n199 < 16; n199 = n199 + 1) 
        begin: outbit199
            assign data_11[n199 + d199*16 + c7*28*16] = data_11_array[c7][d199][n199];
        end
    endgenerate
    generate 
        localparam integer d200 = 4;
        for (n200 = 0; n200 < 16; n200 = n200 + 1) 
        begin: outbit200
            assign data_11[n200 + d200*16 + c7*28*16] = data_11_array[c7][d200][n200];
        end
    endgenerate
    generate 
        localparam integer d201 = 5;
        for (n201 = 0; n201 < 16; n201 = n201 + 1) 
        begin: outbit201
            assign data_11[n201 + d201*16 + c7*28*16] = data_11_array[c7][d201][n201];
        end
    endgenerate
    generate 
        localparam integer d202 = 6;
        for (n202 = 0; n202 < 16; n202 = n202 + 1) 
        begin: outbit202
            assign data_11[n202 + d202*16 + c7*28*16] = data_11_array[c7][d202][n202];
        end
    endgenerate
    generate 
        localparam integer d203 = 7;
        for (n203 = 0; n203 < 16; n203 = n203 + 1) 
        begin: outbit203
            assign data_11[n203 + d203*16 + c7*28*16] = data_11_array[c7][d203][n203];
        end
    endgenerate
    generate 
        localparam integer d204 = 8;
        for (n204 = 0; n204 < 16; n204 = n204 + 1) 
        begin: outbit204
            assign data_11[n204 + d204*16 + c7*28*16] = data_11_array[c7][d204][n204];
        end
    endgenerate
    generate 
        localparam integer d205 = 9;
        for (n205 = 0; n205 < 16; n205 = n205 + 1) 
        begin: outbit205
            assign data_11[n205 + d205*16 + c7*28*16] = data_11_array[c7][d205][n205];
        end
    endgenerate
    generate 
        localparam integer d206 = 10;
        for (n206 = 0; n206 < 16; n206 = n206 + 1) 
        begin: outbit206
            assign data_11[n206 + d206*16 + c7*28*16] = data_11_array[c7][d206][n206];
        end
    endgenerate
    generate 
        localparam integer d207 = 11;
        for (n207 = 0; n207 < 16; n207 = n207 + 1) 
        begin: outbit207
            assign data_11[n207 + d207*16 + c7*28*16] = data_11_array[c7][d207][n207];
        end
    endgenerate
    generate 
        localparam integer d208 = 12;
        for (n208 = 0; n208 < 16; n208 = n208 + 1) 
        begin: outbit208
            assign data_11[n208 + d208*16 + c7*28*16] = data_11_array[c7][d208][n208];
        end
    endgenerate
    generate 
        localparam integer d209 = 13;
        for (n209 = 0; n209 < 16; n209 = n209 + 1) 
        begin: outbit209
            assign data_11[n209 + d209*16 + c7*28*16] = data_11_array[c7][d209][n209];
        end
    endgenerate
    generate 
        localparam integer d210 = 14;
        for (n210 = 0; n210 < 16; n210 = n210 + 1) 
        begin: outbit210
            assign data_11[n210 + d210*16 + c7*28*16] = data_11_array[c7][d210][n210];
        end
    endgenerate
    generate 
        localparam integer d211 = 15;
        for (n211 = 0; n211 < 16; n211 = n211 + 1) 
        begin: outbit211
            assign data_11[n211 + d211*16 + c7*28*16] = data_11_array[c7][d211][n211];
        end
    endgenerate
    generate 
        localparam integer d212 = 16;
        for (n212 = 0; n212 < 16; n212 = n212 + 1) 
        begin: outbit212
            assign data_11[n212 + d212*16 + c7*28*16] = data_11_array[c7][d212][n212];
        end
    endgenerate
    generate 
        localparam integer d213 = 17;
        for (n213 = 0; n213 < 16; n213 = n213 + 1) 
        begin: outbit213
            assign data_11[n213 + d213*16 + c7*28*16] = data_11_array[c7][d213][n213];
        end
    endgenerate
    generate 
        localparam integer d214 = 18;
        for (n214 = 0; n214 < 16; n214 = n214 + 1) 
        begin: outbit214
            assign data_11[n214 + d214*16 + c7*28*16] = data_11_array[c7][d214][n214];
        end
    endgenerate
    generate 
        localparam integer d215 = 19;
        for (n215 = 0; n215 < 16; n215 = n215 + 1) 
        begin: outbit215
            assign data_11[n215 + d215*16 + c7*28*16] = data_11_array[c7][d215][n215];
        end
    endgenerate
    generate 
        localparam integer d216 = 20;
        for (n216 = 0; n216 < 16; n216 = n216 + 1) 
        begin: outbit216
            assign data_11[n216 + d216*16 + c7*28*16] = data_11_array[c7][d216][n216];
        end
    endgenerate
    generate 
        localparam integer d217 = 21;
        for (n217 = 0; n217 < 16; n217 = n217 + 1) 
        begin: outbit217
            assign data_11[n217 + d217*16 + c7*28*16] = data_11_array[c7][d217][n217];
        end
    endgenerate
    generate 
        localparam integer d218 = 22;
        for (n218 = 0; n218 < 16; n218 = n218 + 1) 
        begin: outbit218
            assign data_11[n218 + d218*16 + c7*28*16] = data_11_array[c7][d218][n218];
        end
    endgenerate
    generate 
        localparam integer d219 = 23;
        for (n219 = 0; n219 < 16; n219 = n219 + 1) 
        begin: outbit219
            assign data_11[n219 + d219*16 + c7*28*16] = data_11_array[c7][d219][n219];
        end
    endgenerate
    generate 
        localparam integer d220 = 24;
        for (n220 = 0; n220 < 16; n220 = n220 + 1) 
        begin: outbit220
            assign data_11[n220 + d220*16 + c7*28*16] = data_11_array[c7][d220][n220];
        end
    endgenerate
    generate 
        localparam integer d221 = 25;
        for (n221 = 0; n221 < 16; n221 = n221 + 1) 
        begin: outbit221
            assign data_11[n221 + d221*16 + c7*28*16] = data_11_array[c7][d221][n221];
        end
    endgenerate
    generate 
        localparam integer d222 = 26;
        for (n222 = 0; n222 < 16; n222 = n222 + 1) 
        begin: outbit222
            assign data_11[n222 + d222*16 + c7*28*16] = data_11_array[c7][d222][n222];
        end
    endgenerate
    generate 
        localparam integer d223 = 27;
        for (n223 = 0; n223 < 16; n223 = n223 + 1) 
        begin: outbit223
            assign data_11[n223 + d223*16 + c7*28*16] = data_11_array[c7][d223][n223];
        end
    endgenerate
    localparam integer c8 = 8;
    generate 
        localparam integer d224 = 0;
        for (n224 = 0; n224 < 16; n224 = n224 + 1) 
        begin: outbit224
            assign data_11[n224 + d224*16 + c8*28*16] = data_11_array[c8][d224][n224];
        end
    endgenerate
    generate 
        localparam integer d225 = 1;
        for (n225 = 0; n225 < 16; n225 = n225 + 1) 
        begin: outbit225
            assign data_11[n225 + d225*16 + c8*28*16] = data_11_array[c8][d225][n225];
        end
    endgenerate
    generate 
        localparam integer d226 = 2;
        for (n226 = 0; n226 < 16; n226 = n226 + 1) 
        begin: outbit226
            assign data_11[n226 + d226*16 + c8*28*16] = data_11_array[c8][d226][n226];
        end
    endgenerate
    generate 
        localparam integer d227 = 3;
        for (n227 = 0; n227 < 16; n227 = n227 + 1) 
        begin: outbit227
            assign data_11[n227 + d227*16 + c8*28*16] = data_11_array[c8][d227][n227];
        end
    endgenerate
    generate 
        localparam integer d228 = 4;
        for (n228 = 0; n228 < 16; n228 = n228 + 1) 
        begin: outbit228
            assign data_11[n228 + d228*16 + c8*28*16] = data_11_array[c8][d228][n228];
        end
    endgenerate
    generate 
        localparam integer d229 = 5;
        for (n229 = 0; n229 < 16; n229 = n229 + 1) 
        begin: outbit229
            assign data_11[n229 + d229*16 + c8*28*16] = data_11_array[c8][d229][n229];
        end
    endgenerate
    generate 
        localparam integer d230 = 6;
        for (n230 = 0; n230 < 16; n230 = n230 + 1) 
        begin: outbit230
            assign data_11[n230 + d230*16 + c8*28*16] = data_11_array[c8][d230][n230];
        end
    endgenerate
    generate 
        localparam integer d231 = 7;
        for (n231 = 0; n231 < 16; n231 = n231 + 1) 
        begin: outbit231
            assign data_11[n231 + d231*16 + c8*28*16] = data_11_array[c8][d231][n231];
        end
    endgenerate
    generate 
        localparam integer d232 = 8;
        for (n232 = 0; n232 < 16; n232 = n232 + 1) 
        begin: outbit232
            assign data_11[n232 + d232*16 + c8*28*16] = data_11_array[c8][d232][n232];
        end
    endgenerate
    generate 
        localparam integer d233 = 9;
        for (n233 = 0; n233 < 16; n233 = n233 + 1) 
        begin: outbit233
            assign data_11[n233 + d233*16 + c8*28*16] = data_11_array[c8][d233][n233];
        end
    endgenerate
    generate 
        localparam integer d234 = 10;
        for (n234 = 0; n234 < 16; n234 = n234 + 1) 
        begin: outbit234
            assign data_11[n234 + d234*16 + c8*28*16] = data_11_array[c8][d234][n234];
        end
    endgenerate
    generate 
        localparam integer d235 = 11;
        for (n235 = 0; n235 < 16; n235 = n235 + 1) 
        begin: outbit235
            assign data_11[n235 + d235*16 + c8*28*16] = data_11_array[c8][d235][n235];
        end
    endgenerate
    generate 
        localparam integer d236 = 12;
        for (n236 = 0; n236 < 16; n236 = n236 + 1) 
        begin: outbit236
            assign data_11[n236 + d236*16 + c8*28*16] = data_11_array[c8][d236][n236];
        end
    endgenerate
    generate 
        localparam integer d237 = 13;
        for (n237 = 0; n237 < 16; n237 = n237 + 1) 
        begin: outbit237
            assign data_11[n237 + d237*16 + c8*28*16] = data_11_array[c8][d237][n237];
        end
    endgenerate
    generate 
        localparam integer d238 = 14;
        for (n238 = 0; n238 < 16; n238 = n238 + 1) 
        begin: outbit238
            assign data_11[n238 + d238*16 + c8*28*16] = data_11_array[c8][d238][n238];
        end
    endgenerate
    generate 
        localparam integer d239 = 15;
        for (n239 = 0; n239 < 16; n239 = n239 + 1) 
        begin: outbit239
            assign data_11[n239 + d239*16 + c8*28*16] = data_11_array[c8][d239][n239];
        end
    endgenerate
    generate 
        localparam integer d240 = 16;
        for (n240 = 0; n240 < 16; n240 = n240 + 1) 
        begin: outbit240
            assign data_11[n240 + d240*16 + c8*28*16] = data_11_array[c8][d240][n240];
        end
    endgenerate
    generate 
        localparam integer d241 = 17;
        for (n241 = 0; n241 < 16; n241 = n241 + 1) 
        begin: outbit241
            assign data_11[n241 + d241*16 + c8*28*16] = data_11_array[c8][d241][n241];
        end
    endgenerate
    generate 
        localparam integer d242 = 18;
        for (n242 = 0; n242 < 16; n242 = n242 + 1) 
        begin: outbit242
            assign data_11[n242 + d242*16 + c8*28*16] = data_11_array[c8][d242][n242];
        end
    endgenerate
    generate 
        localparam integer d243 = 19;
        for (n243 = 0; n243 < 16; n243 = n243 + 1) 
        begin: outbit243
            assign data_11[n243 + d243*16 + c8*28*16] = data_11_array[c8][d243][n243];
        end
    endgenerate
    generate 
        localparam integer d244 = 20;
        for (n244 = 0; n244 < 16; n244 = n244 + 1) 
        begin: outbit244
            assign data_11[n244 + d244*16 + c8*28*16] = data_11_array[c8][d244][n244];
        end
    endgenerate
    generate 
        localparam integer d245 = 21;
        for (n245 = 0; n245 < 16; n245 = n245 + 1) 
        begin: outbit245
            assign data_11[n245 + d245*16 + c8*28*16] = data_11_array[c8][d245][n245];
        end
    endgenerate
    generate 
        localparam integer d246 = 22;
        for (n246 = 0; n246 < 16; n246 = n246 + 1) 
        begin: outbit246
            assign data_11[n246 + d246*16 + c8*28*16] = data_11_array[c8][d246][n246];
        end
    endgenerate
    generate 
        localparam integer d247 = 23;
        for (n247 = 0; n247 < 16; n247 = n247 + 1) 
        begin: outbit247
            assign data_11[n247 + d247*16 + c8*28*16] = data_11_array[c8][d247][n247];
        end
    endgenerate
    generate 
        localparam integer d248 = 24;
        for (n248 = 0; n248 < 16; n248 = n248 + 1) 
        begin: outbit248
            assign data_11[n248 + d248*16 + c8*28*16] = data_11_array[c8][d248][n248];
        end
    endgenerate
    generate 
        localparam integer d249 = 25;
        for (n249 = 0; n249 < 16; n249 = n249 + 1) 
        begin: outbit249
            assign data_11[n249 + d249*16 + c8*28*16] = data_11_array[c8][d249][n249];
        end
    endgenerate
    generate 
        localparam integer d250 = 26;
        for (n250 = 0; n250 < 16; n250 = n250 + 1) 
        begin: outbit250
            assign data_11[n250 + d250*16 + c8*28*16] = data_11_array[c8][d250][n250];
        end
    endgenerate
    generate 
        localparam integer d251 = 27;
        for (n251 = 0; n251 < 16; n251 = n251 + 1) 
        begin: outbit251
            assign data_11[n251 + d251*16 + c8*28*16] = data_11_array[c8][d251][n251];
        end
    endgenerate
    localparam integer c9 = 9;
    generate 
        localparam integer d252 = 0;
        for (n252 = 0; n252 < 16; n252 = n252 + 1) 
        begin: outbit252
            assign data_11[n252 + d252*16 + c9*28*16] = data_11_array[c9][d252][n252];
        end
    endgenerate
    generate 
        localparam integer d253 = 1;
        for (n253 = 0; n253 < 16; n253 = n253 + 1) 
        begin: outbit253
            assign data_11[n253 + d253*16 + c9*28*16] = data_11_array[c9][d253][n253];
        end
    endgenerate
    generate 
        localparam integer d254 = 2;
        for (n254 = 0; n254 < 16; n254 = n254 + 1) 
        begin: outbit254
            assign data_11[n254 + d254*16 + c9*28*16] = data_11_array[c9][d254][n254];
        end
    endgenerate
    generate 
        localparam integer d255 = 3;
        for (n255 = 0; n255 < 16; n255 = n255 + 1) 
        begin: outbit255
            assign data_11[n255 + d255*16 + c9*28*16] = data_11_array[c9][d255][n255];
        end
    endgenerate
    generate 
        localparam integer d256 = 4;
        for (n256 = 0; n256 < 16; n256 = n256 + 1) 
        begin: outbit256
            assign data_11[n256 + d256*16 + c9*28*16] = data_11_array[c9][d256][n256];
        end
    endgenerate
    generate 
        localparam integer d257 = 5;
        for (n257 = 0; n257 < 16; n257 = n257 + 1) 
        begin: outbit257
            assign data_11[n257 + d257*16 + c9*28*16] = data_11_array[c9][d257][n257];
        end
    endgenerate
    generate 
        localparam integer d258 = 6;
        for (n258 = 0; n258 < 16; n258 = n258 + 1) 
        begin: outbit258
            assign data_11[n258 + d258*16 + c9*28*16] = data_11_array[c9][d258][n258];
        end
    endgenerate
    generate 
        localparam integer d259 = 7;
        for (n259 = 0; n259 < 16; n259 = n259 + 1) 
        begin: outbit259
            assign data_11[n259 + d259*16 + c9*28*16] = data_11_array[c9][d259][n259];
        end
    endgenerate
    generate 
        localparam integer d260 = 8;
        for (n260 = 0; n260 < 16; n260 = n260 + 1) 
        begin: outbit260
            assign data_11[n260 + d260*16 + c9*28*16] = data_11_array[c9][d260][n260];
        end
    endgenerate
    generate 
        localparam integer d261 = 9;
        for (n261 = 0; n261 < 16; n261 = n261 + 1) 
        begin: outbit261
            assign data_11[n261 + d261*16 + c9*28*16] = data_11_array[c9][d261][n261];
        end
    endgenerate
    generate 
        localparam integer d262 = 10;
        for (n262 = 0; n262 < 16; n262 = n262 + 1) 
        begin: outbit262
            assign data_11[n262 + d262*16 + c9*28*16] = data_11_array[c9][d262][n262];
        end
    endgenerate
    generate 
        localparam integer d263 = 11;
        for (n263 = 0; n263 < 16; n263 = n263 + 1) 
        begin: outbit263
            assign data_11[n263 + d263*16 + c9*28*16] = data_11_array[c9][d263][n263];
        end
    endgenerate
    generate 
        localparam integer d264 = 12;
        for (n264 = 0; n264 < 16; n264 = n264 + 1) 
        begin: outbit264
            assign data_11[n264 + d264*16 + c9*28*16] = data_11_array[c9][d264][n264];
        end
    endgenerate
    generate 
        localparam integer d265 = 13;
        for (n265 = 0; n265 < 16; n265 = n265 + 1) 
        begin: outbit265
            assign data_11[n265 + d265*16 + c9*28*16] = data_11_array[c9][d265][n265];
        end
    endgenerate
    generate 
        localparam integer d266 = 14;
        for (n266 = 0; n266 < 16; n266 = n266 + 1) 
        begin: outbit266
            assign data_11[n266 + d266*16 + c9*28*16] = data_11_array[c9][d266][n266];
        end
    endgenerate
    generate 
        localparam integer d267 = 15;
        for (n267 = 0; n267 < 16; n267 = n267 + 1) 
        begin: outbit267
            assign data_11[n267 + d267*16 + c9*28*16] = data_11_array[c9][d267][n267];
        end
    endgenerate
    generate 
        localparam integer d268 = 16;
        for (n268 = 0; n268 < 16; n268 = n268 + 1) 
        begin: outbit268
            assign data_11[n268 + d268*16 + c9*28*16] = data_11_array[c9][d268][n268];
        end
    endgenerate
    generate 
        localparam integer d269 = 17;
        for (n269 = 0; n269 < 16; n269 = n269 + 1) 
        begin: outbit269
            assign data_11[n269 + d269*16 + c9*28*16] = data_11_array[c9][d269][n269];
        end
    endgenerate
    generate 
        localparam integer d270 = 18;
        for (n270 = 0; n270 < 16; n270 = n270 + 1) 
        begin: outbit270
            assign data_11[n270 + d270*16 + c9*28*16] = data_11_array[c9][d270][n270];
        end
    endgenerate
    generate 
        localparam integer d271 = 19;
        for (n271 = 0; n271 < 16; n271 = n271 + 1) 
        begin: outbit271
            assign data_11[n271 + d271*16 + c9*28*16] = data_11_array[c9][d271][n271];
        end
    endgenerate
    generate 
        localparam integer d272 = 20;
        for (n272 = 0; n272 < 16; n272 = n272 + 1) 
        begin: outbit272
            assign data_11[n272 + d272*16 + c9*28*16] = data_11_array[c9][d272][n272];
        end
    endgenerate
    generate 
        localparam integer d273 = 21;
        for (n273 = 0; n273 < 16; n273 = n273 + 1) 
        begin: outbit273
            assign data_11[n273 + d273*16 + c9*28*16] = data_11_array[c9][d273][n273];
        end
    endgenerate
    generate 
        localparam integer d274 = 22;
        for (n274 = 0; n274 < 16; n274 = n274 + 1) 
        begin: outbit274
            assign data_11[n274 + d274*16 + c9*28*16] = data_11_array[c9][d274][n274];
        end
    endgenerate
    generate 
        localparam integer d275 = 23;
        for (n275 = 0; n275 < 16; n275 = n275 + 1) 
        begin: outbit275
            assign data_11[n275 + d275*16 + c9*28*16] = data_11_array[c9][d275][n275];
        end
    endgenerate
    generate 
        localparam integer d276 = 24;
        for (n276 = 0; n276 < 16; n276 = n276 + 1) 
        begin: outbit276
            assign data_11[n276 + d276*16 + c9*28*16] = data_11_array[c9][d276][n276];
        end
    endgenerate
    generate 
        localparam integer d277 = 25;
        for (n277 = 0; n277 < 16; n277 = n277 + 1) 
        begin: outbit277
            assign data_11[n277 + d277*16 + c9*28*16] = data_11_array[c9][d277][n277];
        end
    endgenerate
    generate 
        localparam integer d278 = 26;
        for (n278 = 0; n278 < 16; n278 = n278 + 1) 
        begin: outbit278
            assign data_11[n278 + d278*16 + c9*28*16] = data_11_array[c9][d278][n278];
        end
    endgenerate
    generate 
        localparam integer d279 = 27;
        for (n279 = 0; n279 < 16; n279 = n279 + 1) 
        begin: outbit279
            assign data_11[n279 + d279*16 + c9*28*16] = data_11_array[c9][d279][n279];
        end
    endgenerate
    localparam integer c10 = 10;
    generate 
        localparam integer d280 = 0;
        for (n280 = 0; n280 < 16; n280 = n280 + 1) 
        begin: outbit280
            assign data_11[n280 + d280*16 + c10*28*16] = data_11_array[c10][d280][n280];
        end
    endgenerate
    generate 
        localparam integer d281 = 1;
        for (n281 = 0; n281 < 16; n281 = n281 + 1) 
        begin: outbit281
            assign data_11[n281 + d281*16 + c10*28*16] = data_11_array[c10][d281][n281];
        end
    endgenerate
    generate 
        localparam integer d282 = 2;
        for (n282 = 0; n282 < 16; n282 = n282 + 1) 
        begin: outbit282
            assign data_11[n282 + d282*16 + c10*28*16] = data_11_array[c10][d282][n282];
        end
    endgenerate
    generate 
        localparam integer d283 = 3;
        for (n283 = 0; n283 < 16; n283 = n283 + 1) 
        begin: outbit283
            assign data_11[n283 + d283*16 + c10*28*16] = data_11_array[c10][d283][n283];
        end
    endgenerate
    generate 
        localparam integer d284 = 4;
        for (n284 = 0; n284 < 16; n284 = n284 + 1) 
        begin: outbit284
            assign data_11[n284 + d284*16 + c10*28*16] = data_11_array[c10][d284][n284];
        end
    endgenerate
    generate 
        localparam integer d285 = 5;
        for (n285 = 0; n285 < 16; n285 = n285 + 1) 
        begin: outbit285
            assign data_11[n285 + d285*16 + c10*28*16] = data_11_array[c10][d285][n285];
        end
    endgenerate
    generate 
        localparam integer d286 = 6;
        for (n286 = 0; n286 < 16; n286 = n286 + 1) 
        begin: outbit286
            assign data_11[n286 + d286*16 + c10*28*16] = data_11_array[c10][d286][n286];
        end
    endgenerate
    generate 
        localparam integer d287 = 7;
        for (n287 = 0; n287 < 16; n287 = n287 + 1) 
        begin: outbit287
            assign data_11[n287 + d287*16 + c10*28*16] = data_11_array[c10][d287][n287];
        end
    endgenerate
    generate 
        localparam integer d288 = 8;
        for (n288 = 0; n288 < 16; n288 = n288 + 1) 
        begin: outbit288
            assign data_11[n288 + d288*16 + c10*28*16] = data_11_array[c10][d288][n288];
        end
    endgenerate
    generate 
        localparam integer d289 = 9;
        for (n289 = 0; n289 < 16; n289 = n289 + 1) 
        begin: outbit289
            assign data_11[n289 + d289*16 + c10*28*16] = data_11_array[c10][d289][n289];
        end
    endgenerate
    generate 
        localparam integer d290 = 10;
        for (n290 = 0; n290 < 16; n290 = n290 + 1) 
        begin: outbit290
            assign data_11[n290 + d290*16 + c10*28*16] = data_11_array[c10][d290][n290];
        end
    endgenerate
    generate 
        localparam integer d291 = 11;
        for (n291 = 0; n291 < 16; n291 = n291 + 1) 
        begin: outbit291
            assign data_11[n291 + d291*16 + c10*28*16] = data_11_array[c10][d291][n291];
        end
    endgenerate
    generate 
        localparam integer d292 = 12;
        for (n292 = 0; n292 < 16; n292 = n292 + 1) 
        begin: outbit292
            assign data_11[n292 + d292*16 + c10*28*16] = data_11_array[c10][d292][n292];
        end
    endgenerate
    generate 
        localparam integer d293 = 13;
        for (n293 = 0; n293 < 16; n293 = n293 + 1) 
        begin: outbit293
            assign data_11[n293 + d293*16 + c10*28*16] = data_11_array[c10][d293][n293];
        end
    endgenerate
    generate 
        localparam integer d294 = 14;
        for (n294 = 0; n294 < 16; n294 = n294 + 1) 
        begin: outbit294
            assign data_11[n294 + d294*16 + c10*28*16] = data_11_array[c10][d294][n294];
        end
    endgenerate
    generate 
        localparam integer d295 = 15;
        for (n295 = 0; n295 < 16; n295 = n295 + 1) 
        begin: outbit295
            assign data_11[n295 + d295*16 + c10*28*16] = data_11_array[c10][d295][n295];
        end
    endgenerate
    generate 
        localparam integer d296 = 16;
        for (n296 = 0; n296 < 16; n296 = n296 + 1) 
        begin: outbit296
            assign data_11[n296 + d296*16 + c10*28*16] = data_11_array[c10][d296][n296];
        end
    endgenerate
    generate 
        localparam integer d297 = 17;
        for (n297 = 0; n297 < 16; n297 = n297 + 1) 
        begin: outbit297
            assign data_11[n297 + d297*16 + c10*28*16] = data_11_array[c10][d297][n297];
        end
    endgenerate
    generate 
        localparam integer d298 = 18;
        for (n298 = 0; n298 < 16; n298 = n298 + 1) 
        begin: outbit298
            assign data_11[n298 + d298*16 + c10*28*16] = data_11_array[c10][d298][n298];
        end
    endgenerate
    generate 
        localparam integer d299 = 19;
        for (n299 = 0; n299 < 16; n299 = n299 + 1) 
        begin: outbit299
            assign data_11[n299 + d299*16 + c10*28*16] = data_11_array[c10][d299][n299];
        end
    endgenerate
    generate 
        localparam integer d300 = 20;
        for (n300 = 0; n300 < 16; n300 = n300 + 1) 
        begin: outbit300
            assign data_11[n300 + d300*16 + c10*28*16] = data_11_array[c10][d300][n300];
        end
    endgenerate
    generate 
        localparam integer d301 = 21;
        for (n301 = 0; n301 < 16; n301 = n301 + 1) 
        begin: outbit301
            assign data_11[n301 + d301*16 + c10*28*16] = data_11_array[c10][d301][n301];
        end
    endgenerate
    generate 
        localparam integer d302 = 22;
        for (n302 = 0; n302 < 16; n302 = n302 + 1) 
        begin: outbit302
            assign data_11[n302 + d302*16 + c10*28*16] = data_11_array[c10][d302][n302];
        end
    endgenerate
    generate 
        localparam integer d303 = 23;
        for (n303 = 0; n303 < 16; n303 = n303 + 1) 
        begin: outbit303
            assign data_11[n303 + d303*16 + c10*28*16] = data_11_array[c10][d303][n303];
        end
    endgenerate
    generate 
        localparam integer d304 = 24;
        for (n304 = 0; n304 < 16; n304 = n304 + 1) 
        begin: outbit304
            assign data_11[n304 + d304*16 + c10*28*16] = data_11_array[c10][d304][n304];
        end
    endgenerate
    generate 
        localparam integer d305 = 25;
        for (n305 = 0; n305 < 16; n305 = n305 + 1) 
        begin: outbit305
            assign data_11[n305 + d305*16 + c10*28*16] = data_11_array[c10][d305][n305];
        end
    endgenerate
    generate 
        localparam integer d306 = 26;
        for (n306 = 0; n306 < 16; n306 = n306 + 1) 
        begin: outbit306
            assign data_11[n306 + d306*16 + c10*28*16] = data_11_array[c10][d306][n306];
        end
    endgenerate
    generate 
        localparam integer d307 = 27;
        for (n307 = 0; n307 < 16; n307 = n307 + 1) 
        begin: outbit307
            assign data_11[n307 + d307*16 + c10*28*16] = data_11_array[c10][d307][n307];
        end
    endgenerate
    localparam integer c11 = 11;
    generate 
        localparam integer d308 = 0;
        for (n308 = 0; n308 < 16; n308 = n308 + 1) 
        begin: outbit308
            assign data_11[n308 + d308*16 + c11*28*16] = data_11_array[c11][d308][n308];
        end
    endgenerate
    generate 
        localparam integer d309 = 1;
        for (n309 = 0; n309 < 16; n309 = n309 + 1) 
        begin: outbit309
            assign data_11[n309 + d309*16 + c11*28*16] = data_11_array[c11][d309][n309];
        end
    endgenerate
    generate 
        localparam integer d310 = 2;
        for (n310 = 0; n310 < 16; n310 = n310 + 1) 
        begin: outbit310
            assign data_11[n310 + d310*16 + c11*28*16] = data_11_array[c11][d310][n310];
        end
    endgenerate
    generate 
        localparam integer d311 = 3;
        for (n311 = 0; n311 < 16; n311 = n311 + 1) 
        begin: outbit311
            assign data_11[n311 + d311*16 + c11*28*16] = data_11_array[c11][d311][n311];
        end
    endgenerate
    generate 
        localparam integer d312 = 4;
        for (n312 = 0; n312 < 16; n312 = n312 + 1) 
        begin: outbit312
            assign data_11[n312 + d312*16 + c11*28*16] = data_11_array[c11][d312][n312];
        end
    endgenerate
    generate 
        localparam integer d313 = 5;
        for (n313 = 0; n313 < 16; n313 = n313 + 1) 
        begin: outbit313
            assign data_11[n313 + d313*16 + c11*28*16] = data_11_array[c11][d313][n313];
        end
    endgenerate
    generate 
        localparam integer d314 = 6;
        for (n314 = 0; n314 < 16; n314 = n314 + 1) 
        begin: outbit314
            assign data_11[n314 + d314*16 + c11*28*16] = data_11_array[c11][d314][n314];
        end
    endgenerate
    generate 
        localparam integer d315 = 7;
        for (n315 = 0; n315 < 16; n315 = n315 + 1) 
        begin: outbit315
            assign data_11[n315 + d315*16 + c11*28*16] = data_11_array[c11][d315][n315];
        end
    endgenerate
    generate 
        localparam integer d316 = 8;
        for (n316 = 0; n316 < 16; n316 = n316 + 1) 
        begin: outbit316
            assign data_11[n316 + d316*16 + c11*28*16] = data_11_array[c11][d316][n316];
        end
    endgenerate
    generate 
        localparam integer d317 = 9;
        for (n317 = 0; n317 < 16; n317 = n317 + 1) 
        begin: outbit317
            assign data_11[n317 + d317*16 + c11*28*16] = data_11_array[c11][d317][n317];
        end
    endgenerate
    generate 
        localparam integer d318 = 10;
        for (n318 = 0; n318 < 16; n318 = n318 + 1) 
        begin: outbit318
            assign data_11[n318 + d318*16 + c11*28*16] = data_11_array[c11][d318][n318];
        end
    endgenerate
    generate 
        localparam integer d319 = 11;
        for (n319 = 0; n319 < 16; n319 = n319 + 1) 
        begin: outbit319
            assign data_11[n319 + d319*16 + c11*28*16] = data_11_array[c11][d319][n319];
        end
    endgenerate
    generate 
        localparam integer d320 = 12;
        for (n320 = 0; n320 < 16; n320 = n320 + 1) 
        begin: outbit320
            assign data_11[n320 + d320*16 + c11*28*16] = data_11_array[c11][d320][n320];
        end
    endgenerate
    generate 
        localparam integer d321 = 13;
        for (n321 = 0; n321 < 16; n321 = n321 + 1) 
        begin: outbit321
            assign data_11[n321 + d321*16 + c11*28*16] = data_11_array[c11][d321][n321];
        end
    endgenerate
    generate 
        localparam integer d322 = 14;
        for (n322 = 0; n322 < 16; n322 = n322 + 1) 
        begin: outbit322
            assign data_11[n322 + d322*16 + c11*28*16] = data_11_array[c11][d322][n322];
        end
    endgenerate
    generate 
        localparam integer d323 = 15;
        for (n323 = 0; n323 < 16; n323 = n323 + 1) 
        begin: outbit323
            assign data_11[n323 + d323*16 + c11*28*16] = data_11_array[c11][d323][n323];
        end
    endgenerate
    generate 
        localparam integer d324 = 16;
        for (n324 = 0; n324 < 16; n324 = n324 + 1) 
        begin: outbit324
            assign data_11[n324 + d324*16 + c11*28*16] = data_11_array[c11][d324][n324];
        end
    endgenerate
    generate 
        localparam integer d325 = 17;
        for (n325 = 0; n325 < 16; n325 = n325 + 1) 
        begin: outbit325
            assign data_11[n325 + d325*16 + c11*28*16] = data_11_array[c11][d325][n325];
        end
    endgenerate
    generate 
        localparam integer d326 = 18;
        for (n326 = 0; n326 < 16; n326 = n326 + 1) 
        begin: outbit326
            assign data_11[n326 + d326*16 + c11*28*16] = data_11_array[c11][d326][n326];
        end
    endgenerate
    generate 
        localparam integer d327 = 19;
        for (n327 = 0; n327 < 16; n327 = n327 + 1) 
        begin: outbit327
            assign data_11[n327 + d327*16 + c11*28*16] = data_11_array[c11][d327][n327];
        end
    endgenerate
    generate 
        localparam integer d328 = 20;
        for (n328 = 0; n328 < 16; n328 = n328 + 1) 
        begin: outbit328
            assign data_11[n328 + d328*16 + c11*28*16] = data_11_array[c11][d328][n328];
        end
    endgenerate
    generate 
        localparam integer d329 = 21;
        for (n329 = 0; n329 < 16; n329 = n329 + 1) 
        begin: outbit329
            assign data_11[n329 + d329*16 + c11*28*16] = data_11_array[c11][d329][n329];
        end
    endgenerate
    generate 
        localparam integer d330 = 22;
        for (n330 = 0; n330 < 16; n330 = n330 + 1) 
        begin: outbit330
            assign data_11[n330 + d330*16 + c11*28*16] = data_11_array[c11][d330][n330];
        end
    endgenerate
    generate 
        localparam integer d331 = 23;
        for (n331 = 0; n331 < 16; n331 = n331 + 1) 
        begin: outbit331
            assign data_11[n331 + d331*16 + c11*28*16] = data_11_array[c11][d331][n331];
        end
    endgenerate
    generate 
        localparam integer d332 = 24;
        for (n332 = 0; n332 < 16; n332 = n332 + 1) 
        begin: outbit332
            assign data_11[n332 + d332*16 + c11*28*16] = data_11_array[c11][d332][n332];
        end
    endgenerate
    generate 
        localparam integer d333 = 25;
        for (n333 = 0; n333 < 16; n333 = n333 + 1) 
        begin: outbit333
            assign data_11[n333 + d333*16 + c11*28*16] = data_11_array[c11][d333][n333];
        end
    endgenerate
    generate 
        localparam integer d334 = 26;
        for (n334 = 0; n334 < 16; n334 = n334 + 1) 
        begin: outbit334
            assign data_11[n334 + d334*16 + c11*28*16] = data_11_array[c11][d334][n334];
        end
    endgenerate
    generate 
        localparam integer d335 = 27;
        for (n335 = 0; n335 < 16; n335 = n335 + 1) 
        begin: outbit335
            assign data_11[n335 + d335*16 + c11*28*16] = data_11_array[c11][d335][n335];
        end
    endgenerate
    localparam integer c12 = 12;
    generate 
        localparam integer d336 = 0;
        for (n336 = 0; n336 < 16; n336 = n336 + 1) 
        begin: outbit336
            assign data_11[n336 + d336*16 + c12*28*16] = data_11_array[c12][d336][n336];
        end
    endgenerate
    generate 
        localparam integer d337 = 1;
        for (n337 = 0; n337 < 16; n337 = n337 + 1) 
        begin: outbit337
            assign data_11[n337 + d337*16 + c12*28*16] = data_11_array[c12][d337][n337];
        end
    endgenerate
    generate 
        localparam integer d338 = 2;
        for (n338 = 0; n338 < 16; n338 = n338 + 1) 
        begin: outbit338
            assign data_11[n338 + d338*16 + c12*28*16] = data_11_array[c12][d338][n338];
        end
    endgenerate
    generate 
        localparam integer d339 = 3;
        for (n339 = 0; n339 < 16; n339 = n339 + 1) 
        begin: outbit339
            assign data_11[n339 + d339*16 + c12*28*16] = data_11_array[c12][d339][n339];
        end
    endgenerate
    generate 
        localparam integer d340 = 4;
        for (n340 = 0; n340 < 16; n340 = n340 + 1) 
        begin: outbit340
            assign data_11[n340 + d340*16 + c12*28*16] = data_11_array[c12][d340][n340];
        end
    endgenerate
    generate 
        localparam integer d341 = 5;
        for (n341 = 0; n341 < 16; n341 = n341 + 1) 
        begin: outbit341
            assign data_11[n341 + d341*16 + c12*28*16] = data_11_array[c12][d341][n341];
        end
    endgenerate
    generate 
        localparam integer d342 = 6;
        for (n342 = 0; n342 < 16; n342 = n342 + 1) 
        begin: outbit342
            assign data_11[n342 + d342*16 + c12*28*16] = data_11_array[c12][d342][n342];
        end
    endgenerate
    generate 
        localparam integer d343 = 7;
        for (n343 = 0; n343 < 16; n343 = n343 + 1) 
        begin: outbit343
            assign data_11[n343 + d343*16 + c12*28*16] = data_11_array[c12][d343][n343];
        end
    endgenerate
    generate 
        localparam integer d344 = 8;
        for (n344 = 0; n344 < 16; n344 = n344 + 1) 
        begin: outbit344
            assign data_11[n344 + d344*16 + c12*28*16] = data_11_array[c12][d344][n344];
        end
    endgenerate
    generate 
        localparam integer d345 = 9;
        for (n345 = 0; n345 < 16; n345 = n345 + 1) 
        begin: outbit345
            assign data_11[n345 + d345*16 + c12*28*16] = data_11_array[c12][d345][n345];
        end
    endgenerate
    generate 
        localparam integer d346 = 10;
        for (n346 = 0; n346 < 16; n346 = n346 + 1) 
        begin: outbit346
            assign data_11[n346 + d346*16 + c12*28*16] = data_11_array[c12][d346][n346];
        end
    endgenerate
    generate 
        localparam integer d347 = 11;
        for (n347 = 0; n347 < 16; n347 = n347 + 1) 
        begin: outbit347
            assign data_11[n347 + d347*16 + c12*28*16] = data_11_array[c12][d347][n347];
        end
    endgenerate
    generate 
        localparam integer d348 = 12;
        for (n348 = 0; n348 < 16; n348 = n348 + 1) 
        begin: outbit348
            assign data_11[n348 + d348*16 + c12*28*16] = data_11_array[c12][d348][n348];
        end
    endgenerate
    generate 
        localparam integer d349 = 13;
        for (n349 = 0; n349 < 16; n349 = n349 + 1) 
        begin: outbit349
            assign data_11[n349 + d349*16 + c12*28*16] = data_11_array[c12][d349][n349];
        end
    endgenerate
    generate 
        localparam integer d350 = 14;
        for (n350 = 0; n350 < 16; n350 = n350 + 1) 
        begin: outbit350
            assign data_11[n350 + d350*16 + c12*28*16] = data_11_array[c12][d350][n350];
        end
    endgenerate
    generate 
        localparam integer d351 = 15;
        for (n351 = 0; n351 < 16; n351 = n351 + 1) 
        begin: outbit351
            assign data_11[n351 + d351*16 + c12*28*16] = data_11_array[c12][d351][n351];
        end
    endgenerate
    generate 
        localparam integer d352 = 16;
        for (n352 = 0; n352 < 16; n352 = n352 + 1) 
        begin: outbit352
            assign data_11[n352 + d352*16 + c12*28*16] = data_11_array[c12][d352][n352];
        end
    endgenerate
    generate 
        localparam integer d353 = 17;
        for (n353 = 0; n353 < 16; n353 = n353 + 1) 
        begin: outbit353
            assign data_11[n353 + d353*16 + c12*28*16] = data_11_array[c12][d353][n353];
        end
    endgenerate
    generate 
        localparam integer d354 = 18;
        for (n354 = 0; n354 < 16; n354 = n354 + 1) 
        begin: outbit354
            assign data_11[n354 + d354*16 + c12*28*16] = data_11_array[c12][d354][n354];
        end
    endgenerate
    generate 
        localparam integer d355 = 19;
        for (n355 = 0; n355 < 16; n355 = n355 + 1) 
        begin: outbit355
            assign data_11[n355 + d355*16 + c12*28*16] = data_11_array[c12][d355][n355];
        end
    endgenerate
    generate 
        localparam integer d356 = 20;
        for (n356 = 0; n356 < 16; n356 = n356 + 1) 
        begin: outbit356
            assign data_11[n356 + d356*16 + c12*28*16] = data_11_array[c12][d356][n356];
        end
    endgenerate
    generate 
        localparam integer d357 = 21;
        for (n357 = 0; n357 < 16; n357 = n357 + 1) 
        begin: outbit357
            assign data_11[n357 + d357*16 + c12*28*16] = data_11_array[c12][d357][n357];
        end
    endgenerate
    generate 
        localparam integer d358 = 22;
        for (n358 = 0; n358 < 16; n358 = n358 + 1) 
        begin: outbit358
            assign data_11[n358 + d358*16 + c12*28*16] = data_11_array[c12][d358][n358];
        end
    endgenerate
    generate 
        localparam integer d359 = 23;
        for (n359 = 0; n359 < 16; n359 = n359 + 1) 
        begin: outbit359
            assign data_11[n359 + d359*16 + c12*28*16] = data_11_array[c12][d359][n359];
        end
    endgenerate
    generate 
        localparam integer d360 = 24;
        for (n360 = 0; n360 < 16; n360 = n360 + 1) 
        begin: outbit360
            assign data_11[n360 + d360*16 + c12*28*16] = data_11_array[c12][d360][n360];
        end
    endgenerate
    generate 
        localparam integer d361 = 25;
        for (n361 = 0; n361 < 16; n361 = n361 + 1) 
        begin: outbit361
            assign data_11[n361 + d361*16 + c12*28*16] = data_11_array[c12][d361][n361];
        end
    endgenerate
    generate 
        localparam integer d362 = 26;
        for (n362 = 0; n362 < 16; n362 = n362 + 1) 
        begin: outbit362
            assign data_11[n362 + d362*16 + c12*28*16] = data_11_array[c12][d362][n362];
        end
    endgenerate
    generate 
        localparam integer d363 = 27;
        for (n363 = 0; n363 < 16; n363 = n363 + 1) 
        begin: outbit363
            assign data_11[n363 + d363*16 + c12*28*16] = data_11_array[c12][d363][n363];
        end
    endgenerate
    localparam integer c13 = 13;
    generate 
        localparam integer d364 = 0;
        for (n364 = 0; n364 < 16; n364 = n364 + 1) 
        begin: outbit364
            assign data_11[n364 + d364*16 + c13*28*16] = data_11_array[c13][d364][n364];
        end
    endgenerate
    generate 
        localparam integer d365 = 1;
        for (n365 = 0; n365 < 16; n365 = n365 + 1) 
        begin: outbit365
            assign data_11[n365 + d365*16 + c13*28*16] = data_11_array[c13][d365][n365];
        end
    endgenerate
    generate 
        localparam integer d366 = 2;
        for (n366 = 0; n366 < 16; n366 = n366 + 1) 
        begin: outbit366
            assign data_11[n366 + d366*16 + c13*28*16] = data_11_array[c13][d366][n366];
        end
    endgenerate
    generate 
        localparam integer d367 = 3;
        for (n367 = 0; n367 < 16; n367 = n367 + 1) 
        begin: outbit367
            assign data_11[n367 + d367*16 + c13*28*16] = data_11_array[c13][d367][n367];
        end
    endgenerate
    generate 
        localparam integer d368 = 4;
        for (n368 = 0; n368 < 16; n368 = n368 + 1) 
        begin: outbit368
            assign data_11[n368 + d368*16 + c13*28*16] = data_11_array[c13][d368][n368];
        end
    endgenerate
    generate 
        localparam integer d369 = 5;
        for (n369 = 0; n369 < 16; n369 = n369 + 1) 
        begin: outbit369
            assign data_11[n369 + d369*16 + c13*28*16] = data_11_array[c13][d369][n369];
        end
    endgenerate
    generate 
        localparam integer d370 = 6;
        for (n370 = 0; n370 < 16; n370 = n370 + 1) 
        begin: outbit370
            assign data_11[n370 + d370*16 + c13*28*16] = data_11_array[c13][d370][n370];
        end
    endgenerate
    generate 
        localparam integer d371 = 7;
        for (n371 = 0; n371 < 16; n371 = n371 + 1) 
        begin: outbit371
            assign data_11[n371 + d371*16 + c13*28*16] = data_11_array[c13][d371][n371];
        end
    endgenerate
    generate 
        localparam integer d372 = 8;
        for (n372 = 0; n372 < 16; n372 = n372 + 1) 
        begin: outbit372
            assign data_11[n372 + d372*16 + c13*28*16] = data_11_array[c13][d372][n372];
        end
    endgenerate
    generate 
        localparam integer d373 = 9;
        for (n373 = 0; n373 < 16; n373 = n373 + 1) 
        begin: outbit373
            assign data_11[n373 + d373*16 + c13*28*16] = data_11_array[c13][d373][n373];
        end
    endgenerate
    generate 
        localparam integer d374 = 10;
        for (n374 = 0; n374 < 16; n374 = n374 + 1) 
        begin: outbit374
            assign data_11[n374 + d374*16 + c13*28*16] = data_11_array[c13][d374][n374];
        end
    endgenerate
    generate 
        localparam integer d375 = 11;
        for (n375 = 0; n375 < 16; n375 = n375 + 1) 
        begin: outbit375
            assign data_11[n375 + d375*16 + c13*28*16] = data_11_array[c13][d375][n375];
        end
    endgenerate
    generate 
        localparam integer d376 = 12;
        for (n376 = 0; n376 < 16; n376 = n376 + 1) 
        begin: outbit376
            assign data_11[n376 + d376*16 + c13*28*16] = data_11_array[c13][d376][n376];
        end
    endgenerate
    generate 
        localparam integer d377 = 13;
        for (n377 = 0; n377 < 16; n377 = n377 + 1) 
        begin: outbit377
            assign data_11[n377 + d377*16 + c13*28*16] = data_11_array[c13][d377][n377];
        end
    endgenerate
    generate 
        localparam integer d378 = 14;
        for (n378 = 0; n378 < 16; n378 = n378 + 1) 
        begin: outbit378
            assign data_11[n378 + d378*16 + c13*28*16] = data_11_array[c13][d378][n378];
        end
    endgenerate
    generate 
        localparam integer d379 = 15;
        for (n379 = 0; n379 < 16; n379 = n379 + 1) 
        begin: outbit379
            assign data_11[n379 + d379*16 + c13*28*16] = data_11_array[c13][d379][n379];
        end
    endgenerate
    generate 
        localparam integer d380 = 16;
        for (n380 = 0; n380 < 16; n380 = n380 + 1) 
        begin: outbit380
            assign data_11[n380 + d380*16 + c13*28*16] = data_11_array[c13][d380][n380];
        end
    endgenerate
    generate 
        localparam integer d381 = 17;
        for (n381 = 0; n381 < 16; n381 = n381 + 1) 
        begin: outbit381
            assign data_11[n381 + d381*16 + c13*28*16] = data_11_array[c13][d381][n381];
        end
    endgenerate
    generate 
        localparam integer d382 = 18;
        for (n382 = 0; n382 < 16; n382 = n382 + 1) 
        begin: outbit382
            assign data_11[n382 + d382*16 + c13*28*16] = data_11_array[c13][d382][n382];
        end
    endgenerate
    generate 
        localparam integer d383 = 19;
        for (n383 = 0; n383 < 16; n383 = n383 + 1) 
        begin: outbit383
            assign data_11[n383 + d383*16 + c13*28*16] = data_11_array[c13][d383][n383];
        end
    endgenerate
    generate 
        localparam integer d384 = 20;
        for (n384 = 0; n384 < 16; n384 = n384 + 1) 
        begin: outbit384
            assign data_11[n384 + d384*16 + c13*28*16] = data_11_array[c13][d384][n384];
        end
    endgenerate
    generate 
        localparam integer d385 = 21;
        for (n385 = 0; n385 < 16; n385 = n385 + 1) 
        begin: outbit385
            assign data_11[n385 + d385*16 + c13*28*16] = data_11_array[c13][d385][n385];
        end
    endgenerate
    generate 
        localparam integer d386 = 22;
        for (n386 = 0; n386 < 16; n386 = n386 + 1) 
        begin: outbit386
            assign data_11[n386 + d386*16 + c13*28*16] = data_11_array[c13][d386][n386];
        end
    endgenerate
    generate 
        localparam integer d387 = 23;
        for (n387 = 0; n387 < 16; n387 = n387 + 1) 
        begin: outbit387
            assign data_11[n387 + d387*16 + c13*28*16] = data_11_array[c13][d387][n387];
        end
    endgenerate
    generate 
        localparam integer d388 = 24;
        for (n388 = 0; n388 < 16; n388 = n388 + 1) 
        begin: outbit388
            assign data_11[n388 + d388*16 + c13*28*16] = data_11_array[c13][d388][n388];
        end
    endgenerate
    generate 
        localparam integer d389 = 25;
        for (n389 = 0; n389 < 16; n389 = n389 + 1) 
        begin: outbit389
            assign data_11[n389 + d389*16 + c13*28*16] = data_11_array[c13][d389][n389];
        end
    endgenerate
    generate 
        localparam integer d390 = 26;
        for (n390 = 0; n390 < 16; n390 = n390 + 1) 
        begin: outbit390
            assign data_11[n390 + d390*16 + c13*28*16] = data_11_array[c13][d390][n390];
        end
    endgenerate
    generate 
        localparam integer d391 = 27;
        for (n391 = 0; n391 < 16; n391 = n391 + 1) 
        begin: outbit391
            assign data_11[n391 + d391*16 + c13*28*16] = data_11_array[c13][d391][n391];
        end
    endgenerate
    localparam integer c14 = 14;
    generate 
        localparam integer d392 = 0;
        for (n392 = 0; n392 < 16; n392 = n392 + 1) 
        begin: outbit392
            assign data_11[n392 + d392*16 + c14*28*16] = data_11_array[c14][d392][n392];
        end
    endgenerate
    generate 
        localparam integer d393 = 1;
        for (n393 = 0; n393 < 16; n393 = n393 + 1) 
        begin: outbit393
            assign data_11[n393 + d393*16 + c14*28*16] = data_11_array[c14][d393][n393];
        end
    endgenerate
    generate 
        localparam integer d394 = 2;
        for (n394 = 0; n394 < 16; n394 = n394 + 1) 
        begin: outbit394
            assign data_11[n394 + d394*16 + c14*28*16] = data_11_array[c14][d394][n394];
        end
    endgenerate
    generate 
        localparam integer d395 = 3;
        for (n395 = 0; n395 < 16; n395 = n395 + 1) 
        begin: outbit395
            assign data_11[n395 + d395*16 + c14*28*16] = data_11_array[c14][d395][n395];
        end
    endgenerate
    generate 
        localparam integer d396 = 4;
        for (n396 = 0; n396 < 16; n396 = n396 + 1) 
        begin: outbit396
            assign data_11[n396 + d396*16 + c14*28*16] = data_11_array[c14][d396][n396];
        end
    endgenerate
    generate 
        localparam integer d397 = 5;
        for (n397 = 0; n397 < 16; n397 = n397 + 1) 
        begin: outbit397
            assign data_11[n397 + d397*16 + c14*28*16] = data_11_array[c14][d397][n397];
        end
    endgenerate
    generate 
        localparam integer d398 = 6;
        for (n398 = 0; n398 < 16; n398 = n398 + 1) 
        begin: outbit398
            assign data_11[n398 + d398*16 + c14*28*16] = data_11_array[c14][d398][n398];
        end
    endgenerate
    generate 
        localparam integer d399 = 7;
        for (n399 = 0; n399 < 16; n399 = n399 + 1) 
        begin: outbit399
            assign data_11[n399 + d399*16 + c14*28*16] = data_11_array[c14][d399][n399];
        end
    endgenerate
    generate 
        localparam integer d400 = 8;
        for (n400 = 0; n400 < 16; n400 = n400 + 1) 
        begin: outbit400
            assign data_11[n400 + d400*16 + c14*28*16] = data_11_array[c14][d400][n400];
        end
    endgenerate
    generate 
        localparam integer d401 = 9;
        for (n401 = 0; n401 < 16; n401 = n401 + 1) 
        begin: outbit401
            assign data_11[n401 + d401*16 + c14*28*16] = data_11_array[c14][d401][n401];
        end
    endgenerate
    generate 
        localparam integer d402 = 10;
        for (n402 = 0; n402 < 16; n402 = n402 + 1) 
        begin: outbit402
            assign data_11[n402 + d402*16 + c14*28*16] = data_11_array[c14][d402][n402];
        end
    endgenerate
    generate 
        localparam integer d403 = 11;
        for (n403 = 0; n403 < 16; n403 = n403 + 1) 
        begin: outbit403
            assign data_11[n403 + d403*16 + c14*28*16] = data_11_array[c14][d403][n403];
        end
    endgenerate
    generate 
        localparam integer d404 = 12;
        for (n404 = 0; n404 < 16; n404 = n404 + 1) 
        begin: outbit404
            assign data_11[n404 + d404*16 + c14*28*16] = data_11_array[c14][d404][n404];
        end
    endgenerate
    generate 
        localparam integer d405 = 13;
        for (n405 = 0; n405 < 16; n405 = n405 + 1) 
        begin: outbit405
            assign data_11[n405 + d405*16 + c14*28*16] = data_11_array[c14][d405][n405];
        end
    endgenerate
    generate 
        localparam integer d406 = 14;
        for (n406 = 0; n406 < 16; n406 = n406 + 1) 
        begin: outbit406
            assign data_11[n406 + d406*16 + c14*28*16] = data_11_array[c14][d406][n406];
        end
    endgenerate
    generate 
        localparam integer d407 = 15;
        for (n407 = 0; n407 < 16; n407 = n407 + 1) 
        begin: outbit407
            assign data_11[n407 + d407*16 + c14*28*16] = data_11_array[c14][d407][n407];
        end
    endgenerate
    generate 
        localparam integer d408 = 16;
        for (n408 = 0; n408 < 16; n408 = n408 + 1) 
        begin: outbit408
            assign data_11[n408 + d408*16 + c14*28*16] = data_11_array[c14][d408][n408];
        end
    endgenerate
    generate 
        localparam integer d409 = 17;
        for (n409 = 0; n409 < 16; n409 = n409 + 1) 
        begin: outbit409
            assign data_11[n409 + d409*16 + c14*28*16] = data_11_array[c14][d409][n409];
        end
    endgenerate
    generate 
        localparam integer d410 = 18;
        for (n410 = 0; n410 < 16; n410 = n410 + 1) 
        begin: outbit410
            assign data_11[n410 + d410*16 + c14*28*16] = data_11_array[c14][d410][n410];
        end
    endgenerate
    generate 
        localparam integer d411 = 19;
        for (n411 = 0; n411 < 16; n411 = n411 + 1) 
        begin: outbit411
            assign data_11[n411 + d411*16 + c14*28*16] = data_11_array[c14][d411][n411];
        end
    endgenerate
    generate 
        localparam integer d412 = 20;
        for (n412 = 0; n412 < 16; n412 = n412 + 1) 
        begin: outbit412
            assign data_11[n412 + d412*16 + c14*28*16] = data_11_array[c14][d412][n412];
        end
    endgenerate
    generate 
        localparam integer d413 = 21;
        for (n413 = 0; n413 < 16; n413 = n413 + 1) 
        begin: outbit413
            assign data_11[n413 + d413*16 + c14*28*16] = data_11_array[c14][d413][n413];
        end
    endgenerate
    generate 
        localparam integer d414 = 22;
        for (n414 = 0; n414 < 16; n414 = n414 + 1) 
        begin: outbit414
            assign data_11[n414 + d414*16 + c14*28*16] = data_11_array[c14][d414][n414];
        end
    endgenerate
    generate 
        localparam integer d415 = 23;
        for (n415 = 0; n415 < 16; n415 = n415 + 1) 
        begin: outbit415
            assign data_11[n415 + d415*16 + c14*28*16] = data_11_array[c14][d415][n415];
        end
    endgenerate
    generate 
        localparam integer d416 = 24;
        for (n416 = 0; n416 < 16; n416 = n416 + 1) 
        begin: outbit416
            assign data_11[n416 + d416*16 + c14*28*16] = data_11_array[c14][d416][n416];
        end
    endgenerate
    generate 
        localparam integer d417 = 25;
        for (n417 = 0; n417 < 16; n417 = n417 + 1) 
        begin: outbit417
            assign data_11[n417 + d417*16 + c14*28*16] = data_11_array[c14][d417][n417];
        end
    endgenerate
    generate 
        localparam integer d418 = 26;
        for (n418 = 0; n418 < 16; n418 = n418 + 1) 
        begin: outbit418
            assign data_11[n418 + d418*16 + c14*28*16] = data_11_array[c14][d418][n418];
        end
    endgenerate
    generate 
        localparam integer d419 = 27;
        for (n419 = 0; n419 < 16; n419 = n419 + 1) 
        begin: outbit419
            assign data_11[n419 + d419*16 + c14*28*16] = data_11_array[c14][d419][n419];
        end
    endgenerate
    localparam integer c15 = 15;
    generate 
        localparam integer d420 = 0;
        for (n420 = 0; n420 < 16; n420 = n420 + 1) 
        begin: outbit420
            assign data_11[n420 + d420*16 + c15*28*16] = data_11_array[c15][d420][n420];
        end
    endgenerate
    generate 
        localparam integer d421 = 1;
        for (n421 = 0; n421 < 16; n421 = n421 + 1) 
        begin: outbit421
            assign data_11[n421 + d421*16 + c15*28*16] = data_11_array[c15][d421][n421];
        end
    endgenerate
    generate 
        localparam integer d422 = 2;
        for (n422 = 0; n422 < 16; n422 = n422 + 1) 
        begin: outbit422
            assign data_11[n422 + d422*16 + c15*28*16] = data_11_array[c15][d422][n422];
        end
    endgenerate
    generate 
        localparam integer d423 = 3;
        for (n423 = 0; n423 < 16; n423 = n423 + 1) 
        begin: outbit423
            assign data_11[n423 + d423*16 + c15*28*16] = data_11_array[c15][d423][n423];
        end
    endgenerate
    generate 
        localparam integer d424 = 4;
        for (n424 = 0; n424 < 16; n424 = n424 + 1) 
        begin: outbit424
            assign data_11[n424 + d424*16 + c15*28*16] = data_11_array[c15][d424][n424];
        end
    endgenerate
    generate 
        localparam integer d425 = 5;
        for (n425 = 0; n425 < 16; n425 = n425 + 1) 
        begin: outbit425
            assign data_11[n425 + d425*16 + c15*28*16] = data_11_array[c15][d425][n425];
        end
    endgenerate
    generate 
        localparam integer d426 = 6;
        for (n426 = 0; n426 < 16; n426 = n426 + 1) 
        begin: outbit426
            assign data_11[n426 + d426*16 + c15*28*16] = data_11_array[c15][d426][n426];
        end
    endgenerate
    generate 
        localparam integer d427 = 7;
        for (n427 = 0; n427 < 16; n427 = n427 + 1) 
        begin: outbit427
            assign data_11[n427 + d427*16 + c15*28*16] = data_11_array[c15][d427][n427];
        end
    endgenerate
    generate 
        localparam integer d428 = 8;
        for (n428 = 0; n428 < 16; n428 = n428 + 1) 
        begin: outbit428
            assign data_11[n428 + d428*16 + c15*28*16] = data_11_array[c15][d428][n428];
        end
    endgenerate
    generate 
        localparam integer d429 = 9;
        for (n429 = 0; n429 < 16; n429 = n429 + 1) 
        begin: outbit429
            assign data_11[n429 + d429*16 + c15*28*16] = data_11_array[c15][d429][n429];
        end
    endgenerate
    generate 
        localparam integer d430 = 10;
        for (n430 = 0; n430 < 16; n430 = n430 + 1) 
        begin: outbit430
            assign data_11[n430 + d430*16 + c15*28*16] = data_11_array[c15][d430][n430];
        end
    endgenerate
    generate 
        localparam integer d431 = 11;
        for (n431 = 0; n431 < 16; n431 = n431 + 1) 
        begin: outbit431
            assign data_11[n431 + d431*16 + c15*28*16] = data_11_array[c15][d431][n431];
        end
    endgenerate
    generate 
        localparam integer d432 = 12;
        for (n432 = 0; n432 < 16; n432 = n432 + 1) 
        begin: outbit432
            assign data_11[n432 + d432*16 + c15*28*16] = data_11_array[c15][d432][n432];
        end
    endgenerate
    generate 
        localparam integer d433 = 13;
        for (n433 = 0; n433 < 16; n433 = n433 + 1) 
        begin: outbit433
            assign data_11[n433 + d433*16 + c15*28*16] = data_11_array[c15][d433][n433];
        end
    endgenerate
    generate 
        localparam integer d434 = 14;
        for (n434 = 0; n434 < 16; n434 = n434 + 1) 
        begin: outbit434
            assign data_11[n434 + d434*16 + c15*28*16] = data_11_array[c15][d434][n434];
        end
    endgenerate
    generate 
        localparam integer d435 = 15;
        for (n435 = 0; n435 < 16; n435 = n435 + 1) 
        begin: outbit435
            assign data_11[n435 + d435*16 + c15*28*16] = data_11_array[c15][d435][n435];
        end
    endgenerate
    generate 
        localparam integer d436 = 16;
        for (n436 = 0; n436 < 16; n436 = n436 + 1) 
        begin: outbit436
            assign data_11[n436 + d436*16 + c15*28*16] = data_11_array[c15][d436][n436];
        end
    endgenerate
    generate 
        localparam integer d437 = 17;
        for (n437 = 0; n437 < 16; n437 = n437 + 1) 
        begin: outbit437
            assign data_11[n437 + d437*16 + c15*28*16] = data_11_array[c15][d437][n437];
        end
    endgenerate
    generate 
        localparam integer d438 = 18;
        for (n438 = 0; n438 < 16; n438 = n438 + 1) 
        begin: outbit438
            assign data_11[n438 + d438*16 + c15*28*16] = data_11_array[c15][d438][n438];
        end
    endgenerate
    generate 
        localparam integer d439 = 19;
        for (n439 = 0; n439 < 16; n439 = n439 + 1) 
        begin: outbit439
            assign data_11[n439 + d439*16 + c15*28*16] = data_11_array[c15][d439][n439];
        end
    endgenerate
    generate 
        localparam integer d440 = 20;
        for (n440 = 0; n440 < 16; n440 = n440 + 1) 
        begin: outbit440
            assign data_11[n440 + d440*16 + c15*28*16] = data_11_array[c15][d440][n440];
        end
    endgenerate
    generate 
        localparam integer d441 = 21;
        for (n441 = 0; n441 < 16; n441 = n441 + 1) 
        begin: outbit441
            assign data_11[n441 + d441*16 + c15*28*16] = data_11_array[c15][d441][n441];
        end
    endgenerate
    generate 
        localparam integer d442 = 22;
        for (n442 = 0; n442 < 16; n442 = n442 + 1) 
        begin: outbit442
            assign data_11[n442 + d442*16 + c15*28*16] = data_11_array[c15][d442][n442];
        end
    endgenerate
    generate 
        localparam integer d443 = 23;
        for (n443 = 0; n443 < 16; n443 = n443 + 1) 
        begin: outbit443
            assign data_11[n443 + d443*16 + c15*28*16] = data_11_array[c15][d443][n443];
        end
    endgenerate
    generate 
        localparam integer d444 = 24;
        for (n444 = 0; n444 < 16; n444 = n444 + 1) 
        begin: outbit444
            assign data_11[n444 + d444*16 + c15*28*16] = data_11_array[c15][d444][n444];
        end
    endgenerate
    generate 
        localparam integer d445 = 25;
        for (n445 = 0; n445 < 16; n445 = n445 + 1) 
        begin: outbit445
            assign data_11[n445 + d445*16 + c15*28*16] = data_11_array[c15][d445][n445];
        end
    endgenerate
    generate 
        localparam integer d446 = 26;
        for (n446 = 0; n446 < 16; n446 = n446 + 1) 
        begin: outbit446
            assign data_11[n446 + d446*16 + c15*28*16] = data_11_array[c15][d446][n446];
        end
    endgenerate
    generate 
        localparam integer d447 = 27;
        for (n447 = 0; n447 < 16; n447 = n447 + 1) 
        begin: outbit447
            assign data_11[n447 + d447*16 + c15*28*16] = data_11_array[c15][d447][n447];
        end
    endgenerate
    localparam integer c16 = 16;
    generate 
        localparam integer d448 = 0;
        for (n448 = 0; n448 < 16; n448 = n448 + 1) 
        begin: outbit448
            assign data_11[n448 + d448*16 + c16*28*16] = data_11_array[c16][d448][n448];
        end
    endgenerate
    generate 
        localparam integer d449 = 1;
        for (n449 = 0; n449 < 16; n449 = n449 + 1) 
        begin: outbit449
            assign data_11[n449 + d449*16 + c16*28*16] = data_11_array[c16][d449][n449];
        end
    endgenerate
    generate 
        localparam integer d450 = 2;
        for (n450 = 0; n450 < 16; n450 = n450 + 1) 
        begin: outbit450
            assign data_11[n450 + d450*16 + c16*28*16] = data_11_array[c16][d450][n450];
        end
    endgenerate
    generate 
        localparam integer d451 = 3;
        for (n451 = 0; n451 < 16; n451 = n451 + 1) 
        begin: outbit451
            assign data_11[n451 + d451*16 + c16*28*16] = data_11_array[c16][d451][n451];
        end
    endgenerate
    generate 
        localparam integer d452 = 4;
        for (n452 = 0; n452 < 16; n452 = n452 + 1) 
        begin: outbit452
            assign data_11[n452 + d452*16 + c16*28*16] = data_11_array[c16][d452][n452];
        end
    endgenerate
    generate 
        localparam integer d453 = 5;
        for (n453 = 0; n453 < 16; n453 = n453 + 1) 
        begin: outbit453
            assign data_11[n453 + d453*16 + c16*28*16] = data_11_array[c16][d453][n453];
        end
    endgenerate
    generate 
        localparam integer d454 = 6;
        for (n454 = 0; n454 < 16; n454 = n454 + 1) 
        begin: outbit454
            assign data_11[n454 + d454*16 + c16*28*16] = data_11_array[c16][d454][n454];
        end
    endgenerate
    generate 
        localparam integer d455 = 7;
        for (n455 = 0; n455 < 16; n455 = n455 + 1) 
        begin: outbit455
            assign data_11[n455 + d455*16 + c16*28*16] = data_11_array[c16][d455][n455];
        end
    endgenerate
    generate 
        localparam integer d456 = 8;
        for (n456 = 0; n456 < 16; n456 = n456 + 1) 
        begin: outbit456
            assign data_11[n456 + d456*16 + c16*28*16] = data_11_array[c16][d456][n456];
        end
    endgenerate
    generate 
        localparam integer d457 = 9;
        for (n457 = 0; n457 < 16; n457 = n457 + 1) 
        begin: outbit457
            assign data_11[n457 + d457*16 + c16*28*16] = data_11_array[c16][d457][n457];
        end
    endgenerate
    generate 
        localparam integer d458 = 10;
        for (n458 = 0; n458 < 16; n458 = n458 + 1) 
        begin: outbit458
            assign data_11[n458 + d458*16 + c16*28*16] = data_11_array[c16][d458][n458];
        end
    endgenerate
    generate 
        localparam integer d459 = 11;
        for (n459 = 0; n459 < 16; n459 = n459 + 1) 
        begin: outbit459
            assign data_11[n459 + d459*16 + c16*28*16] = data_11_array[c16][d459][n459];
        end
    endgenerate
    generate 
        localparam integer d460 = 12;
        for (n460 = 0; n460 < 16; n460 = n460 + 1) 
        begin: outbit460
            assign data_11[n460 + d460*16 + c16*28*16] = data_11_array[c16][d460][n460];
        end
    endgenerate
    generate 
        localparam integer d461 = 13;
        for (n461 = 0; n461 < 16; n461 = n461 + 1) 
        begin: outbit461
            assign data_11[n461 + d461*16 + c16*28*16] = data_11_array[c16][d461][n461];
        end
    endgenerate
    generate 
        localparam integer d462 = 14;
        for (n462 = 0; n462 < 16; n462 = n462 + 1) 
        begin: outbit462
            assign data_11[n462 + d462*16 + c16*28*16] = data_11_array[c16][d462][n462];
        end
    endgenerate
    generate 
        localparam integer d463 = 15;
        for (n463 = 0; n463 < 16; n463 = n463 + 1) 
        begin: outbit463
            assign data_11[n463 + d463*16 + c16*28*16] = data_11_array[c16][d463][n463];
        end
    endgenerate
    generate 
        localparam integer d464 = 16;
        for (n464 = 0; n464 < 16; n464 = n464 + 1) 
        begin: outbit464
            assign data_11[n464 + d464*16 + c16*28*16] = data_11_array[c16][d464][n464];
        end
    endgenerate
    generate 
        localparam integer d465 = 17;
        for (n465 = 0; n465 < 16; n465 = n465 + 1) 
        begin: outbit465
            assign data_11[n465 + d465*16 + c16*28*16] = data_11_array[c16][d465][n465];
        end
    endgenerate
    generate 
        localparam integer d466 = 18;
        for (n466 = 0; n466 < 16; n466 = n466 + 1) 
        begin: outbit466
            assign data_11[n466 + d466*16 + c16*28*16] = data_11_array[c16][d466][n466];
        end
    endgenerate
    generate 
        localparam integer d467 = 19;
        for (n467 = 0; n467 < 16; n467 = n467 + 1) 
        begin: outbit467
            assign data_11[n467 + d467*16 + c16*28*16] = data_11_array[c16][d467][n467];
        end
    endgenerate
    generate 
        localparam integer d468 = 20;
        for (n468 = 0; n468 < 16; n468 = n468 + 1) 
        begin: outbit468
            assign data_11[n468 + d468*16 + c16*28*16] = data_11_array[c16][d468][n468];
        end
    endgenerate
    generate 
        localparam integer d469 = 21;
        for (n469 = 0; n469 < 16; n469 = n469 + 1) 
        begin: outbit469
            assign data_11[n469 + d469*16 + c16*28*16] = data_11_array[c16][d469][n469];
        end
    endgenerate
    generate 
        localparam integer d470 = 22;
        for (n470 = 0; n470 < 16; n470 = n470 + 1) 
        begin: outbit470
            assign data_11[n470 + d470*16 + c16*28*16] = data_11_array[c16][d470][n470];
        end
    endgenerate
    generate 
        localparam integer d471 = 23;
        for (n471 = 0; n471 < 16; n471 = n471 + 1) 
        begin: outbit471
            assign data_11[n471 + d471*16 + c16*28*16] = data_11_array[c16][d471][n471];
        end
    endgenerate
    generate 
        localparam integer d472 = 24;
        for (n472 = 0; n472 < 16; n472 = n472 + 1) 
        begin: outbit472
            assign data_11[n472 + d472*16 + c16*28*16] = data_11_array[c16][d472][n472];
        end
    endgenerate
    generate 
        localparam integer d473 = 25;
        for (n473 = 0; n473 < 16; n473 = n473 + 1) 
        begin: outbit473
            assign data_11[n473 + d473*16 + c16*28*16] = data_11_array[c16][d473][n473];
        end
    endgenerate
    generate 
        localparam integer d474 = 26;
        for (n474 = 0; n474 < 16; n474 = n474 + 1) 
        begin: outbit474
            assign data_11[n474 + d474*16 + c16*28*16] = data_11_array[c16][d474][n474];
        end
    endgenerate
    generate 
        localparam integer d475 = 27;
        for (n475 = 0; n475 < 16; n475 = n475 + 1) 
        begin: outbit475
            assign data_11[n475 + d475*16 + c16*28*16] = data_11_array[c16][d475][n475];
        end
    endgenerate
    localparam integer c17 = 17;
    generate 
        localparam integer d476 = 0;
        for (n476 = 0; n476 < 16; n476 = n476 + 1) 
        begin: outbit476
            assign data_11[n476 + d476*16 + c17*28*16] = data_11_array[c17][d476][n476];
        end
    endgenerate
    generate 
        localparam integer d477 = 1;
        for (n477 = 0; n477 < 16; n477 = n477 + 1) 
        begin: outbit477
            assign data_11[n477 + d477*16 + c17*28*16] = data_11_array[c17][d477][n477];
        end
    endgenerate
    generate 
        localparam integer d478 = 2;
        for (n478 = 0; n478 < 16; n478 = n478 + 1) 
        begin: outbit478
            assign data_11[n478 + d478*16 + c17*28*16] = data_11_array[c17][d478][n478];
        end
    endgenerate
    generate 
        localparam integer d479 = 3;
        for (n479 = 0; n479 < 16; n479 = n479 + 1) 
        begin: outbit479
            assign data_11[n479 + d479*16 + c17*28*16] = data_11_array[c17][d479][n479];
        end
    endgenerate
    generate 
        localparam integer d480 = 4;
        for (n480 = 0; n480 < 16; n480 = n480 + 1) 
        begin: outbit480
            assign data_11[n480 + d480*16 + c17*28*16] = data_11_array[c17][d480][n480];
        end
    endgenerate
    generate 
        localparam integer d481 = 5;
        for (n481 = 0; n481 < 16; n481 = n481 + 1) 
        begin: outbit481
            assign data_11[n481 + d481*16 + c17*28*16] = data_11_array[c17][d481][n481];
        end
    endgenerate
    generate 
        localparam integer d482 = 6;
        for (n482 = 0; n482 < 16; n482 = n482 + 1) 
        begin: outbit482
            assign data_11[n482 + d482*16 + c17*28*16] = data_11_array[c17][d482][n482];
        end
    endgenerate
    generate 
        localparam integer d483 = 7;
        for (n483 = 0; n483 < 16; n483 = n483 + 1) 
        begin: outbit483
            assign data_11[n483 + d483*16 + c17*28*16] = data_11_array[c17][d483][n483];
        end
    endgenerate
    generate 
        localparam integer d484 = 8;
        for (n484 = 0; n484 < 16; n484 = n484 + 1) 
        begin: outbit484
            assign data_11[n484 + d484*16 + c17*28*16] = data_11_array[c17][d484][n484];
        end
    endgenerate
    generate 
        localparam integer d485 = 9;
        for (n485 = 0; n485 < 16; n485 = n485 + 1) 
        begin: outbit485
            assign data_11[n485 + d485*16 + c17*28*16] = data_11_array[c17][d485][n485];
        end
    endgenerate
    generate 
        localparam integer d486 = 10;
        for (n486 = 0; n486 < 16; n486 = n486 + 1) 
        begin: outbit486
            assign data_11[n486 + d486*16 + c17*28*16] = data_11_array[c17][d486][n486];
        end
    endgenerate
    generate 
        localparam integer d487 = 11;
        for (n487 = 0; n487 < 16; n487 = n487 + 1) 
        begin: outbit487
            assign data_11[n487 + d487*16 + c17*28*16] = data_11_array[c17][d487][n487];
        end
    endgenerate
    generate 
        localparam integer d488 = 12;
        for (n488 = 0; n488 < 16; n488 = n488 + 1) 
        begin: outbit488
            assign data_11[n488 + d488*16 + c17*28*16] = data_11_array[c17][d488][n488];
        end
    endgenerate
    generate 
        localparam integer d489 = 13;
        for (n489 = 0; n489 < 16; n489 = n489 + 1) 
        begin: outbit489
            assign data_11[n489 + d489*16 + c17*28*16] = data_11_array[c17][d489][n489];
        end
    endgenerate
    generate 
        localparam integer d490 = 14;
        for (n490 = 0; n490 < 16; n490 = n490 + 1) 
        begin: outbit490
            assign data_11[n490 + d490*16 + c17*28*16] = data_11_array[c17][d490][n490];
        end
    endgenerate
    generate 
        localparam integer d491 = 15;
        for (n491 = 0; n491 < 16; n491 = n491 + 1) 
        begin: outbit491
            assign data_11[n491 + d491*16 + c17*28*16] = data_11_array[c17][d491][n491];
        end
    endgenerate
    generate 
        localparam integer d492 = 16;
        for (n492 = 0; n492 < 16; n492 = n492 + 1) 
        begin: outbit492
            assign data_11[n492 + d492*16 + c17*28*16] = data_11_array[c17][d492][n492];
        end
    endgenerate
    generate 
        localparam integer d493 = 17;
        for (n493 = 0; n493 < 16; n493 = n493 + 1) 
        begin: outbit493
            assign data_11[n493 + d493*16 + c17*28*16] = data_11_array[c17][d493][n493];
        end
    endgenerate
    generate 
        localparam integer d494 = 18;
        for (n494 = 0; n494 < 16; n494 = n494 + 1) 
        begin: outbit494
            assign data_11[n494 + d494*16 + c17*28*16] = data_11_array[c17][d494][n494];
        end
    endgenerate
    generate 
        localparam integer d495 = 19;
        for (n495 = 0; n495 < 16; n495 = n495 + 1) 
        begin: outbit495
            assign data_11[n495 + d495*16 + c17*28*16] = data_11_array[c17][d495][n495];
        end
    endgenerate
    generate 
        localparam integer d496 = 20;
        for (n496 = 0; n496 < 16; n496 = n496 + 1) 
        begin: outbit496
            assign data_11[n496 + d496*16 + c17*28*16] = data_11_array[c17][d496][n496];
        end
    endgenerate
    generate 
        localparam integer d497 = 21;
        for (n497 = 0; n497 < 16; n497 = n497 + 1) 
        begin: outbit497
            assign data_11[n497 + d497*16 + c17*28*16] = data_11_array[c17][d497][n497];
        end
    endgenerate
    generate 
        localparam integer d498 = 22;
        for (n498 = 0; n498 < 16; n498 = n498 + 1) 
        begin: outbit498
            assign data_11[n498 + d498*16 + c17*28*16] = data_11_array[c17][d498][n498];
        end
    endgenerate
    generate 
        localparam integer d499 = 23;
        for (n499 = 0; n499 < 16; n499 = n499 + 1) 
        begin: outbit499
            assign data_11[n499 + d499*16 + c17*28*16] = data_11_array[c17][d499][n499];
        end
    endgenerate
    generate 
        localparam integer d500 = 24;
        for (n500 = 0; n500 < 16; n500 = n500 + 1) 
        begin: outbit500
            assign data_11[n500 + d500*16 + c17*28*16] = data_11_array[c17][d500][n500];
        end
    endgenerate
    generate 
        localparam integer d501 = 25;
        for (n501 = 0; n501 < 16; n501 = n501 + 1) 
        begin: outbit501
            assign data_11[n501 + d501*16 + c17*28*16] = data_11_array[c17][d501][n501];
        end
    endgenerate
    generate 
        localparam integer d502 = 26;
        for (n502 = 0; n502 < 16; n502 = n502 + 1) 
        begin: outbit502
            assign data_11[n502 + d502*16 + c17*28*16] = data_11_array[c17][d502][n502];
        end
    endgenerate
    generate 
        localparam integer d503 = 27;
        for (n503 = 0; n503 < 16; n503 = n503 + 1) 
        begin: outbit503
            assign data_11[n503 + d503*16 + c17*28*16] = data_11_array[c17][d503][n503];
        end
    endgenerate
    localparam integer c18 = 18;
    generate 
        localparam integer d504 = 0;
        for (n504 = 0; n504 < 16; n504 = n504 + 1) 
        begin: outbit504
            assign data_11[n504 + d504*16 + c18*28*16] = data_11_array[c18][d504][n504];
        end
    endgenerate
    generate 
        localparam integer d505 = 1;
        for (n505 = 0; n505 < 16; n505 = n505 + 1) 
        begin: outbit505
            assign data_11[n505 + d505*16 + c18*28*16] = data_11_array[c18][d505][n505];
        end
    endgenerate
    generate 
        localparam integer d506 = 2;
        for (n506 = 0; n506 < 16; n506 = n506 + 1) 
        begin: outbit506
            assign data_11[n506 + d506*16 + c18*28*16] = data_11_array[c18][d506][n506];
        end
    endgenerate
    generate 
        localparam integer d507 = 3;
        for (n507 = 0; n507 < 16; n507 = n507 + 1) 
        begin: outbit507
            assign data_11[n507 + d507*16 + c18*28*16] = data_11_array[c18][d507][n507];
        end
    endgenerate
    generate 
        localparam integer d508 = 4;
        for (n508 = 0; n508 < 16; n508 = n508 + 1) 
        begin: outbit508
            assign data_11[n508 + d508*16 + c18*28*16] = data_11_array[c18][d508][n508];
        end
    endgenerate
    generate 
        localparam integer d509 = 5;
        for (n509 = 0; n509 < 16; n509 = n509 + 1) 
        begin: outbit509
            assign data_11[n509 + d509*16 + c18*28*16] = data_11_array[c18][d509][n509];
        end
    endgenerate
    generate 
        localparam integer d510 = 6;
        for (n510 = 0; n510 < 16; n510 = n510 + 1) 
        begin: outbit510
            assign data_11[n510 + d510*16 + c18*28*16] = data_11_array[c18][d510][n510];
        end
    endgenerate
    generate 
        localparam integer d511 = 7;
        for (n511 = 0; n511 < 16; n511 = n511 + 1) 
        begin: outbit511
            assign data_11[n511 + d511*16 + c18*28*16] = data_11_array[c18][d511][n511];
        end
    endgenerate
    generate 
        localparam integer d512 = 8;
        for (n512 = 0; n512 < 16; n512 = n512 + 1) 
        begin: outbit512
            assign data_11[n512 + d512*16 + c18*28*16] = data_11_array[c18][d512][n512];
        end
    endgenerate
    generate 
        localparam integer d513 = 9;
        for (n513 = 0; n513 < 16; n513 = n513 + 1) 
        begin: outbit513
            assign data_11[n513 + d513*16 + c18*28*16] = data_11_array[c18][d513][n513];
        end
    endgenerate
    generate 
        localparam integer d514 = 10;
        for (n514 = 0; n514 < 16; n514 = n514 + 1) 
        begin: outbit514
            assign data_11[n514 + d514*16 + c18*28*16] = data_11_array[c18][d514][n514];
        end
    endgenerate
    generate 
        localparam integer d515 = 11;
        for (n515 = 0; n515 < 16; n515 = n515 + 1) 
        begin: outbit515
            assign data_11[n515 + d515*16 + c18*28*16] = data_11_array[c18][d515][n515];
        end
    endgenerate
    generate 
        localparam integer d516 = 12;
        for (n516 = 0; n516 < 16; n516 = n516 + 1) 
        begin: outbit516
            assign data_11[n516 + d516*16 + c18*28*16] = data_11_array[c18][d516][n516];
        end
    endgenerate
    generate 
        localparam integer d517 = 13;
        for (n517 = 0; n517 < 16; n517 = n517 + 1) 
        begin: outbit517
            assign data_11[n517 + d517*16 + c18*28*16] = data_11_array[c18][d517][n517];
        end
    endgenerate
    generate 
        localparam integer d518 = 14;
        for (n518 = 0; n518 < 16; n518 = n518 + 1) 
        begin: outbit518
            assign data_11[n518 + d518*16 + c18*28*16] = data_11_array[c18][d518][n518];
        end
    endgenerate
    generate 
        localparam integer d519 = 15;
        for (n519 = 0; n519 < 16; n519 = n519 + 1) 
        begin: outbit519
            assign data_11[n519 + d519*16 + c18*28*16] = data_11_array[c18][d519][n519];
        end
    endgenerate
    generate 
        localparam integer d520 = 16;
        for (n520 = 0; n520 < 16; n520 = n520 + 1) 
        begin: outbit520
            assign data_11[n520 + d520*16 + c18*28*16] = data_11_array[c18][d520][n520];
        end
    endgenerate
    generate 
        localparam integer d521 = 17;
        for (n521 = 0; n521 < 16; n521 = n521 + 1) 
        begin: outbit521
            assign data_11[n521 + d521*16 + c18*28*16] = data_11_array[c18][d521][n521];
        end
    endgenerate
    generate 
        localparam integer d522 = 18;
        for (n522 = 0; n522 < 16; n522 = n522 + 1) 
        begin: outbit522
            assign data_11[n522 + d522*16 + c18*28*16] = data_11_array[c18][d522][n522];
        end
    endgenerate
    generate 
        localparam integer d523 = 19;
        for (n523 = 0; n523 < 16; n523 = n523 + 1) 
        begin: outbit523
            assign data_11[n523 + d523*16 + c18*28*16] = data_11_array[c18][d523][n523];
        end
    endgenerate
    generate 
        localparam integer d524 = 20;
        for (n524 = 0; n524 < 16; n524 = n524 + 1) 
        begin: outbit524
            assign data_11[n524 + d524*16 + c18*28*16] = data_11_array[c18][d524][n524];
        end
    endgenerate
    generate 
        localparam integer d525 = 21;
        for (n525 = 0; n525 < 16; n525 = n525 + 1) 
        begin: outbit525
            assign data_11[n525 + d525*16 + c18*28*16] = data_11_array[c18][d525][n525];
        end
    endgenerate
    generate 
        localparam integer d526 = 22;
        for (n526 = 0; n526 < 16; n526 = n526 + 1) 
        begin: outbit526
            assign data_11[n526 + d526*16 + c18*28*16] = data_11_array[c18][d526][n526];
        end
    endgenerate
    generate 
        localparam integer d527 = 23;
        for (n527 = 0; n527 < 16; n527 = n527 + 1) 
        begin: outbit527
            assign data_11[n527 + d527*16 + c18*28*16] = data_11_array[c18][d527][n527];
        end
    endgenerate
    generate 
        localparam integer d528 = 24;
        for (n528 = 0; n528 < 16; n528 = n528 + 1) 
        begin: outbit528
            assign data_11[n528 + d528*16 + c18*28*16] = data_11_array[c18][d528][n528];
        end
    endgenerate
    generate 
        localparam integer d529 = 25;
        for (n529 = 0; n529 < 16; n529 = n529 + 1) 
        begin: outbit529
            assign data_11[n529 + d529*16 + c18*28*16] = data_11_array[c18][d529][n529];
        end
    endgenerate
    generate 
        localparam integer d530 = 26;
        for (n530 = 0; n530 < 16; n530 = n530 + 1) 
        begin: outbit530
            assign data_11[n530 + d530*16 + c18*28*16] = data_11_array[c18][d530][n530];
        end
    endgenerate
    generate 
        localparam integer d531 = 27;
        for (n531 = 0; n531 < 16; n531 = n531 + 1) 
        begin: outbit531
            assign data_11[n531 + d531*16 + c18*28*16] = data_11_array[c18][d531][n531];
        end
    endgenerate
    localparam integer c19 = 19;
    generate 
        localparam integer d532 = 0;
        for (n532 = 0; n532 < 16; n532 = n532 + 1) 
        begin: outbit532
            assign data_11[n532 + d532*16 + c19*28*16] = data_11_array[c19][d532][n532];
        end
    endgenerate
    generate 
        localparam integer d533 = 1;
        for (n533 = 0; n533 < 16; n533 = n533 + 1) 
        begin: outbit533
            assign data_11[n533 + d533*16 + c19*28*16] = data_11_array[c19][d533][n533];
        end
    endgenerate
    generate 
        localparam integer d534 = 2;
        for (n534 = 0; n534 < 16; n534 = n534 + 1) 
        begin: outbit534
            assign data_11[n534 + d534*16 + c19*28*16] = data_11_array[c19][d534][n534];
        end
    endgenerate
    generate 
        localparam integer d535 = 3;
        for (n535 = 0; n535 < 16; n535 = n535 + 1) 
        begin: outbit535
            assign data_11[n535 + d535*16 + c19*28*16] = data_11_array[c19][d535][n535];
        end
    endgenerate
    generate 
        localparam integer d536 = 4;
        for (n536 = 0; n536 < 16; n536 = n536 + 1) 
        begin: outbit536
            assign data_11[n536 + d536*16 + c19*28*16] = data_11_array[c19][d536][n536];
        end
    endgenerate
    generate 
        localparam integer d537 = 5;
        for (n537 = 0; n537 < 16; n537 = n537 + 1) 
        begin: outbit537
            assign data_11[n537 + d537*16 + c19*28*16] = data_11_array[c19][d537][n537];
        end
    endgenerate
    generate 
        localparam integer d538 = 6;
        for (n538 = 0; n538 < 16; n538 = n538 + 1) 
        begin: outbit538
            assign data_11[n538 + d538*16 + c19*28*16] = data_11_array[c19][d538][n538];
        end
    endgenerate
    generate 
        localparam integer d539 = 7;
        for (n539 = 0; n539 < 16; n539 = n539 + 1) 
        begin: outbit539
            assign data_11[n539 + d539*16 + c19*28*16] = data_11_array[c19][d539][n539];
        end
    endgenerate
    generate 
        localparam integer d540 = 8;
        for (n540 = 0; n540 < 16; n540 = n540 + 1) 
        begin: outbit540
            assign data_11[n540 + d540*16 + c19*28*16] = data_11_array[c19][d540][n540];
        end
    endgenerate
    generate 
        localparam integer d541 = 9;
        for (n541 = 0; n541 < 16; n541 = n541 + 1) 
        begin: outbit541
            assign data_11[n541 + d541*16 + c19*28*16] = data_11_array[c19][d541][n541];
        end
    endgenerate
    generate 
        localparam integer d542 = 10;
        for (n542 = 0; n542 < 16; n542 = n542 + 1) 
        begin: outbit542
            assign data_11[n542 + d542*16 + c19*28*16] = data_11_array[c19][d542][n542];
        end
    endgenerate
    generate 
        localparam integer d543 = 11;
        for (n543 = 0; n543 < 16; n543 = n543 + 1) 
        begin: outbit543
            assign data_11[n543 + d543*16 + c19*28*16] = data_11_array[c19][d543][n543];
        end
    endgenerate
    generate 
        localparam integer d544 = 12;
        for (n544 = 0; n544 < 16; n544 = n544 + 1) 
        begin: outbit544
            assign data_11[n544 + d544*16 + c19*28*16] = data_11_array[c19][d544][n544];
        end
    endgenerate
    generate 
        localparam integer d545 = 13;
        for (n545 = 0; n545 < 16; n545 = n545 + 1) 
        begin: outbit545
            assign data_11[n545 + d545*16 + c19*28*16] = data_11_array[c19][d545][n545];
        end
    endgenerate
    generate 
        localparam integer d546 = 14;
        for (n546 = 0; n546 < 16; n546 = n546 + 1) 
        begin: outbit546
            assign data_11[n546 + d546*16 + c19*28*16] = data_11_array[c19][d546][n546];
        end
    endgenerate
    generate 
        localparam integer d547 = 15;
        for (n547 = 0; n547 < 16; n547 = n547 + 1) 
        begin: outbit547
            assign data_11[n547 + d547*16 + c19*28*16] = data_11_array[c19][d547][n547];
        end
    endgenerate
    generate 
        localparam integer d548 = 16;
        for (n548 = 0; n548 < 16; n548 = n548 + 1) 
        begin: outbit548
            assign data_11[n548 + d548*16 + c19*28*16] = data_11_array[c19][d548][n548];
        end
    endgenerate
    generate 
        localparam integer d549 = 17;
        for (n549 = 0; n549 < 16; n549 = n549 + 1) 
        begin: outbit549
            assign data_11[n549 + d549*16 + c19*28*16] = data_11_array[c19][d549][n549];
        end
    endgenerate
    generate 
        localparam integer d550 = 18;
        for (n550 = 0; n550 < 16; n550 = n550 + 1) 
        begin: outbit550
            assign data_11[n550 + d550*16 + c19*28*16] = data_11_array[c19][d550][n550];
        end
    endgenerate
    generate 
        localparam integer d551 = 19;
        for (n551 = 0; n551 < 16; n551 = n551 + 1) 
        begin: outbit551
            assign data_11[n551 + d551*16 + c19*28*16] = data_11_array[c19][d551][n551];
        end
    endgenerate
    generate 
        localparam integer d552 = 20;
        for (n552 = 0; n552 < 16; n552 = n552 + 1) 
        begin: outbit552
            assign data_11[n552 + d552*16 + c19*28*16] = data_11_array[c19][d552][n552];
        end
    endgenerate
    generate 
        localparam integer d553 = 21;
        for (n553 = 0; n553 < 16; n553 = n553 + 1) 
        begin: outbit553
            assign data_11[n553 + d553*16 + c19*28*16] = data_11_array[c19][d553][n553];
        end
    endgenerate
    generate 
        localparam integer d554 = 22;
        for (n554 = 0; n554 < 16; n554 = n554 + 1) 
        begin: outbit554
            assign data_11[n554 + d554*16 + c19*28*16] = data_11_array[c19][d554][n554];
        end
    endgenerate
    generate 
        localparam integer d555 = 23;
        for (n555 = 0; n555 < 16; n555 = n555 + 1) 
        begin: outbit555
            assign data_11[n555 + d555*16 + c19*28*16] = data_11_array[c19][d555][n555];
        end
    endgenerate
    generate 
        localparam integer d556 = 24;
        for (n556 = 0; n556 < 16; n556 = n556 + 1) 
        begin: outbit556
            assign data_11[n556 + d556*16 + c19*28*16] = data_11_array[c19][d556][n556];
        end
    endgenerate
    generate 
        localparam integer d557 = 25;
        for (n557 = 0; n557 < 16; n557 = n557 + 1) 
        begin: outbit557
            assign data_11[n557 + d557*16 + c19*28*16] = data_11_array[c19][d557][n557];
        end
    endgenerate
    generate 
        localparam integer d558 = 26;
        for (n558 = 0; n558 < 16; n558 = n558 + 1) 
        begin: outbit558
            assign data_11[n558 + d558*16 + c19*28*16] = data_11_array[c19][d558][n558];
        end
    endgenerate
    generate 
        localparam integer d559 = 27;
        for (n559 = 0; n559 < 16; n559 = n559 + 1) 
        begin: outbit559
            assign data_11[n559 + d559*16 + c19*28*16] = data_11_array[c19][d559][n559];
        end
    endgenerate
    localparam integer c20 = 20;
    generate 
        localparam integer d560 = 0;
        for (n560 = 0; n560 < 16; n560 = n560 + 1) 
        begin: outbit560
            assign data_11[n560 + d560*16 + c20*28*16] = data_11_array[c20][d560][n560];
        end
    endgenerate
    generate 
        localparam integer d561 = 1;
        for (n561 = 0; n561 < 16; n561 = n561 + 1) 
        begin: outbit561
            assign data_11[n561 + d561*16 + c20*28*16] = data_11_array[c20][d561][n561];
        end
    endgenerate
    generate 
        localparam integer d562 = 2;
        for (n562 = 0; n562 < 16; n562 = n562 + 1) 
        begin: outbit562
            assign data_11[n562 + d562*16 + c20*28*16] = data_11_array[c20][d562][n562];
        end
    endgenerate
    generate 
        localparam integer d563 = 3;
        for (n563 = 0; n563 < 16; n563 = n563 + 1) 
        begin: outbit563
            assign data_11[n563 + d563*16 + c20*28*16] = data_11_array[c20][d563][n563];
        end
    endgenerate
    generate 
        localparam integer d564 = 4;
        for (n564 = 0; n564 < 16; n564 = n564 + 1) 
        begin: outbit564
            assign data_11[n564 + d564*16 + c20*28*16] = data_11_array[c20][d564][n564];
        end
    endgenerate
    generate 
        localparam integer d565 = 5;
        for (n565 = 0; n565 < 16; n565 = n565 + 1) 
        begin: outbit565
            assign data_11[n565 + d565*16 + c20*28*16] = data_11_array[c20][d565][n565];
        end
    endgenerate
    generate 
        localparam integer d566 = 6;
        for (n566 = 0; n566 < 16; n566 = n566 + 1) 
        begin: outbit566
            assign data_11[n566 + d566*16 + c20*28*16] = data_11_array[c20][d566][n566];
        end
    endgenerate
    generate 
        localparam integer d567 = 7;
        for (n567 = 0; n567 < 16; n567 = n567 + 1) 
        begin: outbit567
            assign data_11[n567 + d567*16 + c20*28*16] = data_11_array[c20][d567][n567];
        end
    endgenerate
    generate 
        localparam integer d568 = 8;
        for (n568 = 0; n568 < 16; n568 = n568 + 1) 
        begin: outbit568
            assign data_11[n568 + d568*16 + c20*28*16] = data_11_array[c20][d568][n568];
        end
    endgenerate
    generate 
        localparam integer d569 = 9;
        for (n569 = 0; n569 < 16; n569 = n569 + 1) 
        begin: outbit569
            assign data_11[n569 + d569*16 + c20*28*16] = data_11_array[c20][d569][n569];
        end
    endgenerate
    generate 
        localparam integer d570 = 10;
        for (n570 = 0; n570 < 16; n570 = n570 + 1) 
        begin: outbit570
            assign data_11[n570 + d570*16 + c20*28*16] = data_11_array[c20][d570][n570];
        end
    endgenerate
    generate 
        localparam integer d571 = 11;
        for (n571 = 0; n571 < 16; n571 = n571 + 1) 
        begin: outbit571
            assign data_11[n571 + d571*16 + c20*28*16] = data_11_array[c20][d571][n571];
        end
    endgenerate
    generate 
        localparam integer d572 = 12;
        for (n572 = 0; n572 < 16; n572 = n572 + 1) 
        begin: outbit572
            assign data_11[n572 + d572*16 + c20*28*16] = data_11_array[c20][d572][n572];
        end
    endgenerate
    generate 
        localparam integer d573 = 13;
        for (n573 = 0; n573 < 16; n573 = n573 + 1) 
        begin: outbit573
            assign data_11[n573 + d573*16 + c20*28*16] = data_11_array[c20][d573][n573];
        end
    endgenerate
    generate 
        localparam integer d574 = 14;
        for (n574 = 0; n574 < 16; n574 = n574 + 1) 
        begin: outbit574
            assign data_11[n574 + d574*16 + c20*28*16] = data_11_array[c20][d574][n574];
        end
    endgenerate
    generate 
        localparam integer d575 = 15;
        for (n575 = 0; n575 < 16; n575 = n575 + 1) 
        begin: outbit575
            assign data_11[n575 + d575*16 + c20*28*16] = data_11_array[c20][d575][n575];
        end
    endgenerate
    generate 
        localparam integer d576 = 16;
        for (n576 = 0; n576 < 16; n576 = n576 + 1) 
        begin: outbit576
            assign data_11[n576 + d576*16 + c20*28*16] = data_11_array[c20][d576][n576];
        end
    endgenerate
    generate 
        localparam integer d577 = 17;
        for (n577 = 0; n577 < 16; n577 = n577 + 1) 
        begin: outbit577
            assign data_11[n577 + d577*16 + c20*28*16] = data_11_array[c20][d577][n577];
        end
    endgenerate
    generate 
        localparam integer d578 = 18;
        for (n578 = 0; n578 < 16; n578 = n578 + 1) 
        begin: outbit578
            assign data_11[n578 + d578*16 + c20*28*16] = data_11_array[c20][d578][n578];
        end
    endgenerate
    generate 
        localparam integer d579 = 19;
        for (n579 = 0; n579 < 16; n579 = n579 + 1) 
        begin: outbit579
            assign data_11[n579 + d579*16 + c20*28*16] = data_11_array[c20][d579][n579];
        end
    endgenerate
    generate 
        localparam integer d580 = 20;
        for (n580 = 0; n580 < 16; n580 = n580 + 1) 
        begin: outbit580
            assign data_11[n580 + d580*16 + c20*28*16] = data_11_array[c20][d580][n580];
        end
    endgenerate
    generate 
        localparam integer d581 = 21;
        for (n581 = 0; n581 < 16; n581 = n581 + 1) 
        begin: outbit581
            assign data_11[n581 + d581*16 + c20*28*16] = data_11_array[c20][d581][n581];
        end
    endgenerate
    generate 
        localparam integer d582 = 22;
        for (n582 = 0; n582 < 16; n582 = n582 + 1) 
        begin: outbit582
            assign data_11[n582 + d582*16 + c20*28*16] = data_11_array[c20][d582][n582];
        end
    endgenerate
    generate 
        localparam integer d583 = 23;
        for (n583 = 0; n583 < 16; n583 = n583 + 1) 
        begin: outbit583
            assign data_11[n583 + d583*16 + c20*28*16] = data_11_array[c20][d583][n583];
        end
    endgenerate
    generate 
        localparam integer d584 = 24;
        for (n584 = 0; n584 < 16; n584 = n584 + 1) 
        begin: outbit584
            assign data_11[n584 + d584*16 + c20*28*16] = data_11_array[c20][d584][n584];
        end
    endgenerate
    generate 
        localparam integer d585 = 25;
        for (n585 = 0; n585 < 16; n585 = n585 + 1) 
        begin: outbit585
            assign data_11[n585 + d585*16 + c20*28*16] = data_11_array[c20][d585][n585];
        end
    endgenerate
    generate 
        localparam integer d586 = 26;
        for (n586 = 0; n586 < 16; n586 = n586 + 1) 
        begin: outbit586
            assign data_11[n586 + d586*16 + c20*28*16] = data_11_array[c20][d586][n586];
        end
    endgenerate
    generate 
        localparam integer d587 = 27;
        for (n587 = 0; n587 < 16; n587 = n587 + 1) 
        begin: outbit587
            assign data_11[n587 + d587*16 + c20*28*16] = data_11_array[c20][d587][n587];
        end
    endgenerate
    localparam integer c21 = 21;
    generate 
        localparam integer d588 = 0;
        for (n588 = 0; n588 < 16; n588 = n588 + 1) 
        begin: outbit588
            assign data_11[n588 + d588*16 + c21*28*16] = data_11_array[c21][d588][n588];
        end
    endgenerate
    generate 
        localparam integer d589 = 1;
        for (n589 = 0; n589 < 16; n589 = n589 + 1) 
        begin: outbit589
            assign data_11[n589 + d589*16 + c21*28*16] = data_11_array[c21][d589][n589];
        end
    endgenerate
    generate 
        localparam integer d590 = 2;
        for (n590 = 0; n590 < 16; n590 = n590 + 1) 
        begin: outbit590
            assign data_11[n590 + d590*16 + c21*28*16] = data_11_array[c21][d590][n590];
        end
    endgenerate
    generate 
        localparam integer d591 = 3;
        for (n591 = 0; n591 < 16; n591 = n591 + 1) 
        begin: outbit591
            assign data_11[n591 + d591*16 + c21*28*16] = data_11_array[c21][d591][n591];
        end
    endgenerate
    generate 
        localparam integer d592 = 4;
        for (n592 = 0; n592 < 16; n592 = n592 + 1) 
        begin: outbit592
            assign data_11[n592 + d592*16 + c21*28*16] = data_11_array[c21][d592][n592];
        end
    endgenerate
    generate 
        localparam integer d593 = 5;
        for (n593 = 0; n593 < 16; n593 = n593 + 1) 
        begin: outbit593
            assign data_11[n593 + d593*16 + c21*28*16] = data_11_array[c21][d593][n593];
        end
    endgenerate
    generate 
        localparam integer d594 = 6;
        for (n594 = 0; n594 < 16; n594 = n594 + 1) 
        begin: outbit594
            assign data_11[n594 + d594*16 + c21*28*16] = data_11_array[c21][d594][n594];
        end
    endgenerate
    generate 
        localparam integer d595 = 7;
        for (n595 = 0; n595 < 16; n595 = n595 + 1) 
        begin: outbit595
            assign data_11[n595 + d595*16 + c21*28*16] = data_11_array[c21][d595][n595];
        end
    endgenerate
    generate 
        localparam integer d596 = 8;
        for (n596 = 0; n596 < 16; n596 = n596 + 1) 
        begin: outbit596
            assign data_11[n596 + d596*16 + c21*28*16] = data_11_array[c21][d596][n596];
        end
    endgenerate
    generate 
        localparam integer d597 = 9;
        for (n597 = 0; n597 < 16; n597 = n597 + 1) 
        begin: outbit597
            assign data_11[n597 + d597*16 + c21*28*16] = data_11_array[c21][d597][n597];
        end
    endgenerate
    generate 
        localparam integer d598 = 10;
        for (n598 = 0; n598 < 16; n598 = n598 + 1) 
        begin: outbit598
            assign data_11[n598 + d598*16 + c21*28*16] = data_11_array[c21][d598][n598];
        end
    endgenerate
    generate 
        localparam integer d599 = 11;
        for (n599 = 0; n599 < 16; n599 = n599 + 1) 
        begin: outbit599
            assign data_11[n599 + d599*16 + c21*28*16] = data_11_array[c21][d599][n599];
        end
    endgenerate
    generate 
        localparam integer d600 = 12;
        for (n600 = 0; n600 < 16; n600 = n600 + 1) 
        begin: outbit600
            assign data_11[n600 + d600*16 + c21*28*16] = data_11_array[c21][d600][n600];
        end
    endgenerate
    generate 
        localparam integer d601 = 13;
        for (n601 = 0; n601 < 16; n601 = n601 + 1) 
        begin: outbit601
            assign data_11[n601 + d601*16 + c21*28*16] = data_11_array[c21][d601][n601];
        end
    endgenerate
    generate 
        localparam integer d602 = 14;
        for (n602 = 0; n602 < 16; n602 = n602 + 1) 
        begin: outbit602
            assign data_11[n602 + d602*16 + c21*28*16] = data_11_array[c21][d602][n602];
        end
    endgenerate
    generate 
        localparam integer d603 = 15;
        for (n603 = 0; n603 < 16; n603 = n603 + 1) 
        begin: outbit603
            assign data_11[n603 + d603*16 + c21*28*16] = data_11_array[c21][d603][n603];
        end
    endgenerate
    generate 
        localparam integer d604 = 16;
        for (n604 = 0; n604 < 16; n604 = n604 + 1) 
        begin: outbit604
            assign data_11[n604 + d604*16 + c21*28*16] = data_11_array[c21][d604][n604];
        end
    endgenerate
    generate 
        localparam integer d605 = 17;
        for (n605 = 0; n605 < 16; n605 = n605 + 1) 
        begin: outbit605
            assign data_11[n605 + d605*16 + c21*28*16] = data_11_array[c21][d605][n605];
        end
    endgenerate
    generate 
        localparam integer d606 = 18;
        for (n606 = 0; n606 < 16; n606 = n606 + 1) 
        begin: outbit606
            assign data_11[n606 + d606*16 + c21*28*16] = data_11_array[c21][d606][n606];
        end
    endgenerate
    generate 
        localparam integer d607 = 19;
        for (n607 = 0; n607 < 16; n607 = n607 + 1) 
        begin: outbit607
            assign data_11[n607 + d607*16 + c21*28*16] = data_11_array[c21][d607][n607];
        end
    endgenerate
    generate 
        localparam integer d608 = 20;
        for (n608 = 0; n608 < 16; n608 = n608 + 1) 
        begin: outbit608
            assign data_11[n608 + d608*16 + c21*28*16] = data_11_array[c21][d608][n608];
        end
    endgenerate
    generate 
        localparam integer d609 = 21;
        for (n609 = 0; n609 < 16; n609 = n609 + 1) 
        begin: outbit609
            assign data_11[n609 + d609*16 + c21*28*16] = data_11_array[c21][d609][n609];
        end
    endgenerate
    generate 
        localparam integer d610 = 22;
        for (n610 = 0; n610 < 16; n610 = n610 + 1) 
        begin: outbit610
            assign data_11[n610 + d610*16 + c21*28*16] = data_11_array[c21][d610][n610];
        end
    endgenerate
    generate 
        localparam integer d611 = 23;
        for (n611 = 0; n611 < 16; n611 = n611 + 1) 
        begin: outbit611
            assign data_11[n611 + d611*16 + c21*28*16] = data_11_array[c21][d611][n611];
        end
    endgenerate
    generate 
        localparam integer d612 = 24;
        for (n612 = 0; n612 < 16; n612 = n612 + 1) 
        begin: outbit612
            assign data_11[n612 + d612*16 + c21*28*16] = data_11_array[c21][d612][n612];
        end
    endgenerate
    generate 
        localparam integer d613 = 25;
        for (n613 = 0; n613 < 16; n613 = n613 + 1) 
        begin: outbit613
            assign data_11[n613 + d613*16 + c21*28*16] = data_11_array[c21][d613][n613];
        end
    endgenerate
    generate 
        localparam integer d614 = 26;
        for (n614 = 0; n614 < 16; n614 = n614 + 1) 
        begin: outbit614
            assign data_11[n614 + d614*16 + c21*28*16] = data_11_array[c21][d614][n614];
        end
    endgenerate
    generate 
        localparam integer d615 = 27;
        for (n615 = 0; n615 < 16; n615 = n615 + 1) 
        begin: outbit615
            assign data_11[n615 + d615*16 + c21*28*16] = data_11_array[c21][d615][n615];
        end
    endgenerate
    localparam integer c22 = 22;
    generate 
        localparam integer d616 = 0;
        for (n616 = 0; n616 < 16; n616 = n616 + 1) 
        begin: outbit616
            assign data_11[n616 + d616*16 + c22*28*16] = data_11_array[c22][d616][n616];
        end
    endgenerate
    generate 
        localparam integer d617 = 1;
        for (n617 = 0; n617 < 16; n617 = n617 + 1) 
        begin: outbit617
            assign data_11[n617 + d617*16 + c22*28*16] = data_11_array[c22][d617][n617];
        end
    endgenerate
    generate 
        localparam integer d618 = 2;
        for (n618 = 0; n618 < 16; n618 = n618 + 1) 
        begin: outbit618
            assign data_11[n618 + d618*16 + c22*28*16] = data_11_array[c22][d618][n618];
        end
    endgenerate
    generate 
        localparam integer d619 = 3;
        for (n619 = 0; n619 < 16; n619 = n619 + 1) 
        begin: outbit619
            assign data_11[n619 + d619*16 + c22*28*16] = data_11_array[c22][d619][n619];
        end
    endgenerate
    generate 
        localparam integer d620 = 4;
        for (n620 = 0; n620 < 16; n620 = n620 + 1) 
        begin: outbit620
            assign data_11[n620 + d620*16 + c22*28*16] = data_11_array[c22][d620][n620];
        end
    endgenerate
    generate 
        localparam integer d621 = 5;
        for (n621 = 0; n621 < 16; n621 = n621 + 1) 
        begin: outbit621
            assign data_11[n621 + d621*16 + c22*28*16] = data_11_array[c22][d621][n621];
        end
    endgenerate
    generate 
        localparam integer d622 = 6;
        for (n622 = 0; n622 < 16; n622 = n622 + 1) 
        begin: outbit622
            assign data_11[n622 + d622*16 + c22*28*16] = data_11_array[c22][d622][n622];
        end
    endgenerate
    generate 
        localparam integer d623 = 7;
        for (n623 = 0; n623 < 16; n623 = n623 + 1) 
        begin: outbit623
            assign data_11[n623 + d623*16 + c22*28*16] = data_11_array[c22][d623][n623];
        end
    endgenerate
    generate 
        localparam integer d624 = 8;
        for (n624 = 0; n624 < 16; n624 = n624 + 1) 
        begin: outbit624
            assign data_11[n624 + d624*16 + c22*28*16] = data_11_array[c22][d624][n624];
        end
    endgenerate
    generate 
        localparam integer d625 = 9;
        for (n625 = 0; n625 < 16; n625 = n625 + 1) 
        begin: outbit625
            assign data_11[n625 + d625*16 + c22*28*16] = data_11_array[c22][d625][n625];
        end
    endgenerate
    generate 
        localparam integer d626 = 10;
        for (n626 = 0; n626 < 16; n626 = n626 + 1) 
        begin: outbit626
            assign data_11[n626 + d626*16 + c22*28*16] = data_11_array[c22][d626][n626];
        end
    endgenerate
    generate 
        localparam integer d627 = 11;
        for (n627 = 0; n627 < 16; n627 = n627 + 1) 
        begin: outbit627
            assign data_11[n627 + d627*16 + c22*28*16] = data_11_array[c22][d627][n627];
        end
    endgenerate
    generate 
        localparam integer d628 = 12;
        for (n628 = 0; n628 < 16; n628 = n628 + 1) 
        begin: outbit628
            assign data_11[n628 + d628*16 + c22*28*16] = data_11_array[c22][d628][n628];
        end
    endgenerate
    generate 
        localparam integer d629 = 13;
        for (n629 = 0; n629 < 16; n629 = n629 + 1) 
        begin: outbit629
            assign data_11[n629 + d629*16 + c22*28*16] = data_11_array[c22][d629][n629];
        end
    endgenerate
    generate 
        localparam integer d630 = 14;
        for (n630 = 0; n630 < 16; n630 = n630 + 1) 
        begin: outbit630
            assign data_11[n630 + d630*16 + c22*28*16] = data_11_array[c22][d630][n630];
        end
    endgenerate
    generate 
        localparam integer d631 = 15;
        for (n631 = 0; n631 < 16; n631 = n631 + 1) 
        begin: outbit631
            assign data_11[n631 + d631*16 + c22*28*16] = data_11_array[c22][d631][n631];
        end
    endgenerate
    generate 
        localparam integer d632 = 16;
        for (n632 = 0; n632 < 16; n632 = n632 + 1) 
        begin: outbit632
            assign data_11[n632 + d632*16 + c22*28*16] = data_11_array[c22][d632][n632];
        end
    endgenerate
    generate 
        localparam integer d633 = 17;
        for (n633 = 0; n633 < 16; n633 = n633 + 1) 
        begin: outbit633
            assign data_11[n633 + d633*16 + c22*28*16] = data_11_array[c22][d633][n633];
        end
    endgenerate
    generate 
        localparam integer d634 = 18;
        for (n634 = 0; n634 < 16; n634 = n634 + 1) 
        begin: outbit634
            assign data_11[n634 + d634*16 + c22*28*16] = data_11_array[c22][d634][n634];
        end
    endgenerate
    generate 
        localparam integer d635 = 19;
        for (n635 = 0; n635 < 16; n635 = n635 + 1) 
        begin: outbit635
            assign data_11[n635 + d635*16 + c22*28*16] = data_11_array[c22][d635][n635];
        end
    endgenerate
    generate 
        localparam integer d636 = 20;
        for (n636 = 0; n636 < 16; n636 = n636 + 1) 
        begin: outbit636
            assign data_11[n636 + d636*16 + c22*28*16] = data_11_array[c22][d636][n636];
        end
    endgenerate
    generate 
        localparam integer d637 = 21;
        for (n637 = 0; n637 < 16; n637 = n637 + 1) 
        begin: outbit637
            assign data_11[n637 + d637*16 + c22*28*16] = data_11_array[c22][d637][n637];
        end
    endgenerate
    generate 
        localparam integer d638 = 22;
        for (n638 = 0; n638 < 16; n638 = n638 + 1) 
        begin: outbit638
            assign data_11[n638 + d638*16 + c22*28*16] = data_11_array[c22][d638][n638];
        end
    endgenerate
    generate 
        localparam integer d639 = 23;
        for (n639 = 0; n639 < 16; n639 = n639 + 1) 
        begin: outbit639
            assign data_11[n639 + d639*16 + c22*28*16] = data_11_array[c22][d639][n639];
        end
    endgenerate
    generate 
        localparam integer d640 = 24;
        for (n640 = 0; n640 < 16; n640 = n640 + 1) 
        begin: outbit640
            assign data_11[n640 + d640*16 + c22*28*16] = data_11_array[c22][d640][n640];
        end
    endgenerate
    generate 
        localparam integer d641 = 25;
        for (n641 = 0; n641 < 16; n641 = n641 + 1) 
        begin: outbit641
            assign data_11[n641 + d641*16 + c22*28*16] = data_11_array[c22][d641][n641];
        end
    endgenerate
    generate 
        localparam integer d642 = 26;
        for (n642 = 0; n642 < 16; n642 = n642 + 1) 
        begin: outbit642
            assign data_11[n642 + d642*16 + c22*28*16] = data_11_array[c22][d642][n642];
        end
    endgenerate
    generate 
        localparam integer d643 = 27;
        for (n643 = 0; n643 < 16; n643 = n643 + 1) 
        begin: outbit643
            assign data_11[n643 + d643*16 + c22*28*16] = data_11_array[c22][d643][n643];
        end
    endgenerate
    localparam integer c23 = 23;
    generate 
        localparam integer d644 = 0;
        for (n644 = 0; n644 < 16; n644 = n644 + 1) 
        begin: outbit644
            assign data_11[n644 + d644*16 + c23*28*16] = data_11_array[c23][d644][n644];
        end
    endgenerate
    generate 
        localparam integer d645 = 1;
        for (n645 = 0; n645 < 16; n645 = n645 + 1) 
        begin: outbit645
            assign data_11[n645 + d645*16 + c23*28*16] = data_11_array[c23][d645][n645];
        end
    endgenerate
    generate 
        localparam integer d646 = 2;
        for (n646 = 0; n646 < 16; n646 = n646 + 1) 
        begin: outbit646
            assign data_11[n646 + d646*16 + c23*28*16] = data_11_array[c23][d646][n646];
        end
    endgenerate
    generate 
        localparam integer d647 = 3;
        for (n647 = 0; n647 < 16; n647 = n647 + 1) 
        begin: outbit647
            assign data_11[n647 + d647*16 + c23*28*16] = data_11_array[c23][d647][n647];
        end
    endgenerate
    generate 
        localparam integer d648 = 4;
        for (n648 = 0; n648 < 16; n648 = n648 + 1) 
        begin: outbit648
            assign data_11[n648 + d648*16 + c23*28*16] = data_11_array[c23][d648][n648];
        end
    endgenerate
    generate 
        localparam integer d649 = 5;
        for (n649 = 0; n649 < 16; n649 = n649 + 1) 
        begin: outbit649
            assign data_11[n649 + d649*16 + c23*28*16] = data_11_array[c23][d649][n649];
        end
    endgenerate
    generate 
        localparam integer d650 = 6;
        for (n650 = 0; n650 < 16; n650 = n650 + 1) 
        begin: outbit650
            assign data_11[n650 + d650*16 + c23*28*16] = data_11_array[c23][d650][n650];
        end
    endgenerate
    generate 
        localparam integer d651 = 7;
        for (n651 = 0; n651 < 16; n651 = n651 + 1) 
        begin: outbit651
            assign data_11[n651 + d651*16 + c23*28*16] = data_11_array[c23][d651][n651];
        end
    endgenerate
    generate 
        localparam integer d652 = 8;
        for (n652 = 0; n652 < 16; n652 = n652 + 1) 
        begin: outbit652
            assign data_11[n652 + d652*16 + c23*28*16] = data_11_array[c23][d652][n652];
        end
    endgenerate
    generate 
        localparam integer d653 = 9;
        for (n653 = 0; n653 < 16; n653 = n653 + 1) 
        begin: outbit653
            assign data_11[n653 + d653*16 + c23*28*16] = data_11_array[c23][d653][n653];
        end
    endgenerate
    generate 
        localparam integer d654 = 10;
        for (n654 = 0; n654 < 16; n654 = n654 + 1) 
        begin: outbit654
            assign data_11[n654 + d654*16 + c23*28*16] = data_11_array[c23][d654][n654];
        end
    endgenerate
    generate 
        localparam integer d655 = 11;
        for (n655 = 0; n655 < 16; n655 = n655 + 1) 
        begin: outbit655
            assign data_11[n655 + d655*16 + c23*28*16] = data_11_array[c23][d655][n655];
        end
    endgenerate
    generate 
        localparam integer d656 = 12;
        for (n656 = 0; n656 < 16; n656 = n656 + 1) 
        begin: outbit656
            assign data_11[n656 + d656*16 + c23*28*16] = data_11_array[c23][d656][n656];
        end
    endgenerate
    generate 
        localparam integer d657 = 13;
        for (n657 = 0; n657 < 16; n657 = n657 + 1) 
        begin: outbit657
            assign data_11[n657 + d657*16 + c23*28*16] = data_11_array[c23][d657][n657];
        end
    endgenerate
    generate 
        localparam integer d658 = 14;
        for (n658 = 0; n658 < 16; n658 = n658 + 1) 
        begin: outbit658
            assign data_11[n658 + d658*16 + c23*28*16] = data_11_array[c23][d658][n658];
        end
    endgenerate
    generate 
        localparam integer d659 = 15;
        for (n659 = 0; n659 < 16; n659 = n659 + 1) 
        begin: outbit659
            assign data_11[n659 + d659*16 + c23*28*16] = data_11_array[c23][d659][n659];
        end
    endgenerate
    generate 
        localparam integer d660 = 16;
        for (n660 = 0; n660 < 16; n660 = n660 + 1) 
        begin: outbit660
            assign data_11[n660 + d660*16 + c23*28*16] = data_11_array[c23][d660][n660];
        end
    endgenerate
    generate 
        localparam integer d661 = 17;
        for (n661 = 0; n661 < 16; n661 = n661 + 1) 
        begin: outbit661
            assign data_11[n661 + d661*16 + c23*28*16] = data_11_array[c23][d661][n661];
        end
    endgenerate
    generate 
        localparam integer d662 = 18;
        for (n662 = 0; n662 < 16; n662 = n662 + 1) 
        begin: outbit662
            assign data_11[n662 + d662*16 + c23*28*16] = data_11_array[c23][d662][n662];
        end
    endgenerate
    generate 
        localparam integer d663 = 19;
        for (n663 = 0; n663 < 16; n663 = n663 + 1) 
        begin: outbit663
            assign data_11[n663 + d663*16 + c23*28*16] = data_11_array[c23][d663][n663];
        end
    endgenerate
    generate 
        localparam integer d664 = 20;
        for (n664 = 0; n664 < 16; n664 = n664 + 1) 
        begin: outbit664
            assign data_11[n664 + d664*16 + c23*28*16] = data_11_array[c23][d664][n664];
        end
    endgenerate
    generate 
        localparam integer d665 = 21;
        for (n665 = 0; n665 < 16; n665 = n665 + 1) 
        begin: outbit665
            assign data_11[n665 + d665*16 + c23*28*16] = data_11_array[c23][d665][n665];
        end
    endgenerate
    generate 
        localparam integer d666 = 22;
        for (n666 = 0; n666 < 16; n666 = n666 + 1) 
        begin: outbit666
            assign data_11[n666 + d666*16 + c23*28*16] = data_11_array[c23][d666][n666];
        end
    endgenerate
    generate 
        localparam integer d667 = 23;
        for (n667 = 0; n667 < 16; n667 = n667 + 1) 
        begin: outbit667
            assign data_11[n667 + d667*16 + c23*28*16] = data_11_array[c23][d667][n667];
        end
    endgenerate
    generate 
        localparam integer d668 = 24;
        for (n668 = 0; n668 < 16; n668 = n668 + 1) 
        begin: outbit668
            assign data_11[n668 + d668*16 + c23*28*16] = data_11_array[c23][d668][n668];
        end
    endgenerate
    generate 
        localparam integer d669 = 25;
        for (n669 = 0; n669 < 16; n669 = n669 + 1) 
        begin: outbit669
            assign data_11[n669 + d669*16 + c23*28*16] = data_11_array[c23][d669][n669];
        end
    endgenerate
    generate 
        localparam integer d670 = 26;
        for (n670 = 0; n670 < 16; n670 = n670 + 1) 
        begin: outbit670
            assign data_11[n670 + d670*16 + c23*28*16] = data_11_array[c23][d670][n670];
        end
    endgenerate
    generate 
        localparam integer d671 = 27;
        for (n671 = 0; n671 < 16; n671 = n671 + 1) 
        begin: outbit671
            assign data_11[n671 + d671*16 + c23*28*16] = data_11_array[c23][d671][n671];
        end
    endgenerate
    localparam integer c24 = 24;
    generate 
        localparam integer d672 = 0;
        for (n672 = 0; n672 < 16; n672 = n672 + 1) 
        begin: outbit672
            assign data_11[n672 + d672*16 + c24*28*16] = data_11_array[c24][d672][n672];
        end
    endgenerate
    generate 
        localparam integer d673 = 1;
        for (n673 = 0; n673 < 16; n673 = n673 + 1) 
        begin: outbit673
            assign data_11[n673 + d673*16 + c24*28*16] = data_11_array[c24][d673][n673];
        end
    endgenerate
    generate 
        localparam integer d674 = 2;
        for (n674 = 0; n674 < 16; n674 = n674 + 1) 
        begin: outbit674
            assign data_11[n674 + d674*16 + c24*28*16] = data_11_array[c24][d674][n674];
        end
    endgenerate
    generate 
        localparam integer d675 = 3;
        for (n675 = 0; n675 < 16; n675 = n675 + 1) 
        begin: outbit675
            assign data_11[n675 + d675*16 + c24*28*16] = data_11_array[c24][d675][n675];
        end
    endgenerate
    generate 
        localparam integer d676 = 4;
        for (n676 = 0; n676 < 16; n676 = n676 + 1) 
        begin: outbit676
            assign data_11[n676 + d676*16 + c24*28*16] = data_11_array[c24][d676][n676];
        end
    endgenerate
    generate 
        localparam integer d677 = 5;
        for (n677 = 0; n677 < 16; n677 = n677 + 1) 
        begin: outbit677
            assign data_11[n677 + d677*16 + c24*28*16] = data_11_array[c24][d677][n677];
        end
    endgenerate
    generate 
        localparam integer d678 = 6;
        for (n678 = 0; n678 < 16; n678 = n678 + 1) 
        begin: outbit678
            assign data_11[n678 + d678*16 + c24*28*16] = data_11_array[c24][d678][n678];
        end
    endgenerate
    generate 
        localparam integer d679 = 7;
        for (n679 = 0; n679 < 16; n679 = n679 + 1) 
        begin: outbit679
            assign data_11[n679 + d679*16 + c24*28*16] = data_11_array[c24][d679][n679];
        end
    endgenerate
    generate 
        localparam integer d680 = 8;
        for (n680 = 0; n680 < 16; n680 = n680 + 1) 
        begin: outbit680
            assign data_11[n680 + d680*16 + c24*28*16] = data_11_array[c24][d680][n680];
        end
    endgenerate
    generate 
        localparam integer d681 = 9;
        for (n681 = 0; n681 < 16; n681 = n681 + 1) 
        begin: outbit681
            assign data_11[n681 + d681*16 + c24*28*16] = data_11_array[c24][d681][n681];
        end
    endgenerate
    generate 
        localparam integer d682 = 10;
        for (n682 = 0; n682 < 16; n682 = n682 + 1) 
        begin: outbit682
            assign data_11[n682 + d682*16 + c24*28*16] = data_11_array[c24][d682][n682];
        end
    endgenerate
    generate 
        localparam integer d683 = 11;
        for (n683 = 0; n683 < 16; n683 = n683 + 1) 
        begin: outbit683
            assign data_11[n683 + d683*16 + c24*28*16] = data_11_array[c24][d683][n683];
        end
    endgenerate
    generate 
        localparam integer d684 = 12;
        for (n684 = 0; n684 < 16; n684 = n684 + 1) 
        begin: outbit684
            assign data_11[n684 + d684*16 + c24*28*16] = data_11_array[c24][d684][n684];
        end
    endgenerate
    generate 
        localparam integer d685 = 13;
        for (n685 = 0; n685 < 16; n685 = n685 + 1) 
        begin: outbit685
            assign data_11[n685 + d685*16 + c24*28*16] = data_11_array[c24][d685][n685];
        end
    endgenerate
    generate 
        localparam integer d686 = 14;
        for (n686 = 0; n686 < 16; n686 = n686 + 1) 
        begin: outbit686
            assign data_11[n686 + d686*16 + c24*28*16] = data_11_array[c24][d686][n686];
        end
    endgenerate
    generate 
        localparam integer d687 = 15;
        for (n687 = 0; n687 < 16; n687 = n687 + 1) 
        begin: outbit687
            assign data_11[n687 + d687*16 + c24*28*16] = data_11_array[c24][d687][n687];
        end
    endgenerate
    generate 
        localparam integer d688 = 16;
        for (n688 = 0; n688 < 16; n688 = n688 + 1) 
        begin: outbit688
            assign data_11[n688 + d688*16 + c24*28*16] = data_11_array[c24][d688][n688];
        end
    endgenerate
    generate 
        localparam integer d689 = 17;
        for (n689 = 0; n689 < 16; n689 = n689 + 1) 
        begin: outbit689
            assign data_11[n689 + d689*16 + c24*28*16] = data_11_array[c24][d689][n689];
        end
    endgenerate
    generate 
        localparam integer d690 = 18;
        for (n690 = 0; n690 < 16; n690 = n690 + 1) 
        begin: outbit690
            assign data_11[n690 + d690*16 + c24*28*16] = data_11_array[c24][d690][n690];
        end
    endgenerate
    generate 
        localparam integer d691 = 19;
        for (n691 = 0; n691 < 16; n691 = n691 + 1) 
        begin: outbit691
            assign data_11[n691 + d691*16 + c24*28*16] = data_11_array[c24][d691][n691];
        end
    endgenerate
    generate 
        localparam integer d692 = 20;
        for (n692 = 0; n692 < 16; n692 = n692 + 1) 
        begin: outbit692
            assign data_11[n692 + d692*16 + c24*28*16] = data_11_array[c24][d692][n692];
        end
    endgenerate
    generate 
        localparam integer d693 = 21;
        for (n693 = 0; n693 < 16; n693 = n693 + 1) 
        begin: outbit693
            assign data_11[n693 + d693*16 + c24*28*16] = data_11_array[c24][d693][n693];
        end
    endgenerate
    generate 
        localparam integer d694 = 22;
        for (n694 = 0; n694 < 16; n694 = n694 + 1) 
        begin: outbit694
            assign data_11[n694 + d694*16 + c24*28*16] = data_11_array[c24][d694][n694];
        end
    endgenerate
    generate 
        localparam integer d695 = 23;
        for (n695 = 0; n695 < 16; n695 = n695 + 1) 
        begin: outbit695
            assign data_11[n695 + d695*16 + c24*28*16] = data_11_array[c24][d695][n695];
        end
    endgenerate
    generate 
        localparam integer d696 = 24;
        for (n696 = 0; n696 < 16; n696 = n696 + 1) 
        begin: outbit696
            assign data_11[n696 + d696*16 + c24*28*16] = data_11_array[c24][d696][n696];
        end
    endgenerate
    generate 
        localparam integer d697 = 25;
        for (n697 = 0; n697 < 16; n697 = n697 + 1) 
        begin: outbit697
            assign data_11[n697 + d697*16 + c24*28*16] = data_11_array[c24][d697][n697];
        end
    endgenerate
    generate 
        localparam integer d698 = 26;
        for (n698 = 0; n698 < 16; n698 = n698 + 1) 
        begin: outbit698
            assign data_11[n698 + d698*16 + c24*28*16] = data_11_array[c24][d698][n698];
        end
    endgenerate
    generate 
        localparam integer d699 = 27;
        for (n699 = 0; n699 < 16; n699 = n699 + 1) 
        begin: outbit699
            assign data_11[n699 + d699*16 + c24*28*16] = data_11_array[c24][d699][n699];
        end
    endgenerate
    localparam integer c25 = 25;
    generate 
        localparam integer d700 = 0;
        for (n700 = 0; n700 < 16; n700 = n700 + 1) 
        begin: outbit700
            assign data_11[n700 + d700*16 + c25*28*16] = data_11_array[c25][d700][n700];
        end
    endgenerate
    generate 
        localparam integer d701 = 1;
        for (n701 = 0; n701 < 16; n701 = n701 + 1) 
        begin: outbit701
            assign data_11[n701 + d701*16 + c25*28*16] = data_11_array[c25][d701][n701];
        end
    endgenerate
    generate 
        localparam integer d702 = 2;
        for (n702 = 0; n702 < 16; n702 = n702 + 1) 
        begin: outbit702
            assign data_11[n702 + d702*16 + c25*28*16] = data_11_array[c25][d702][n702];
        end
    endgenerate
    generate 
        localparam integer d703 = 3;
        for (n703 = 0; n703 < 16; n703 = n703 + 1) 
        begin: outbit703
            assign data_11[n703 + d703*16 + c25*28*16] = data_11_array[c25][d703][n703];
        end
    endgenerate
    generate 
        localparam integer d704 = 4;
        for (n704 = 0; n704 < 16; n704 = n704 + 1) 
        begin: outbit704
            assign data_11[n704 + d704*16 + c25*28*16] = data_11_array[c25][d704][n704];
        end
    endgenerate
    generate 
        localparam integer d705 = 5;
        for (n705 = 0; n705 < 16; n705 = n705 + 1) 
        begin: outbit705
            assign data_11[n705 + d705*16 + c25*28*16] = data_11_array[c25][d705][n705];
        end
    endgenerate
    generate 
        localparam integer d706 = 6;
        for (n706 = 0; n706 < 16; n706 = n706 + 1) 
        begin: outbit706
            assign data_11[n706 + d706*16 + c25*28*16] = data_11_array[c25][d706][n706];
        end
    endgenerate
    generate 
        localparam integer d707 = 7;
        for (n707 = 0; n707 < 16; n707 = n707 + 1) 
        begin: outbit707
            assign data_11[n707 + d707*16 + c25*28*16] = data_11_array[c25][d707][n707];
        end
    endgenerate
    generate 
        localparam integer d708 = 8;
        for (n708 = 0; n708 < 16; n708 = n708 + 1) 
        begin: outbit708
            assign data_11[n708 + d708*16 + c25*28*16] = data_11_array[c25][d708][n708];
        end
    endgenerate
    generate 
        localparam integer d709 = 9;
        for (n709 = 0; n709 < 16; n709 = n709 + 1) 
        begin: outbit709
            assign data_11[n709 + d709*16 + c25*28*16] = data_11_array[c25][d709][n709];
        end
    endgenerate
    generate 
        localparam integer d710 = 10;
        for (n710 = 0; n710 < 16; n710 = n710 + 1) 
        begin: outbit710
            assign data_11[n710 + d710*16 + c25*28*16] = data_11_array[c25][d710][n710];
        end
    endgenerate
    generate 
        localparam integer d711 = 11;
        for (n711 = 0; n711 < 16; n711 = n711 + 1) 
        begin: outbit711
            assign data_11[n711 + d711*16 + c25*28*16] = data_11_array[c25][d711][n711];
        end
    endgenerate
    generate 
        localparam integer d712 = 12;
        for (n712 = 0; n712 < 16; n712 = n712 + 1) 
        begin: outbit712
            assign data_11[n712 + d712*16 + c25*28*16] = data_11_array[c25][d712][n712];
        end
    endgenerate
    generate 
        localparam integer d713 = 13;
        for (n713 = 0; n713 < 16; n713 = n713 + 1) 
        begin: outbit713
            assign data_11[n713 + d713*16 + c25*28*16] = data_11_array[c25][d713][n713];
        end
    endgenerate
    generate 
        localparam integer d714 = 14;
        for (n714 = 0; n714 < 16; n714 = n714 + 1) 
        begin: outbit714
            assign data_11[n714 + d714*16 + c25*28*16] = data_11_array[c25][d714][n714];
        end
    endgenerate
    generate 
        localparam integer d715 = 15;
        for (n715 = 0; n715 < 16; n715 = n715 + 1) 
        begin: outbit715
            assign data_11[n715 + d715*16 + c25*28*16] = data_11_array[c25][d715][n715];
        end
    endgenerate
    generate 
        localparam integer d716 = 16;
        for (n716 = 0; n716 < 16; n716 = n716 + 1) 
        begin: outbit716
            assign data_11[n716 + d716*16 + c25*28*16] = data_11_array[c25][d716][n716];
        end
    endgenerate
    generate 
        localparam integer d717 = 17;
        for (n717 = 0; n717 < 16; n717 = n717 + 1) 
        begin: outbit717
            assign data_11[n717 + d717*16 + c25*28*16] = data_11_array[c25][d717][n717];
        end
    endgenerate
    generate 
        localparam integer d718 = 18;
        for (n718 = 0; n718 < 16; n718 = n718 + 1) 
        begin: outbit718
            assign data_11[n718 + d718*16 + c25*28*16] = data_11_array[c25][d718][n718];
        end
    endgenerate
    generate 
        localparam integer d719 = 19;
        for (n719 = 0; n719 < 16; n719 = n719 + 1) 
        begin: outbit719
            assign data_11[n719 + d719*16 + c25*28*16] = data_11_array[c25][d719][n719];
        end
    endgenerate
    generate 
        localparam integer d720 = 20;
        for (n720 = 0; n720 < 16; n720 = n720 + 1) 
        begin: outbit720
            assign data_11[n720 + d720*16 + c25*28*16] = data_11_array[c25][d720][n720];
        end
    endgenerate
    generate 
        localparam integer d721 = 21;
        for (n721 = 0; n721 < 16; n721 = n721 + 1) 
        begin: outbit721
            assign data_11[n721 + d721*16 + c25*28*16] = data_11_array[c25][d721][n721];
        end
    endgenerate
    generate 
        localparam integer d722 = 22;
        for (n722 = 0; n722 < 16; n722 = n722 + 1) 
        begin: outbit722
            assign data_11[n722 + d722*16 + c25*28*16] = data_11_array[c25][d722][n722];
        end
    endgenerate
    generate 
        localparam integer d723 = 23;
        for (n723 = 0; n723 < 16; n723 = n723 + 1) 
        begin: outbit723
            assign data_11[n723 + d723*16 + c25*28*16] = data_11_array[c25][d723][n723];
        end
    endgenerate
    generate 
        localparam integer d724 = 24;
        for (n724 = 0; n724 < 16; n724 = n724 + 1) 
        begin: outbit724
            assign data_11[n724 + d724*16 + c25*28*16] = data_11_array[c25][d724][n724];
        end
    endgenerate
    generate 
        localparam integer d725 = 25;
        for (n725 = 0; n725 < 16; n725 = n725 + 1) 
        begin: outbit725
            assign data_11[n725 + d725*16 + c25*28*16] = data_11_array[c25][d725][n725];
        end
    endgenerate
    generate 
        localparam integer d726 = 26;
        for (n726 = 0; n726 < 16; n726 = n726 + 1) 
        begin: outbit726
            assign data_11[n726 + d726*16 + c25*28*16] = data_11_array[c25][d726][n726];
        end
    endgenerate
    generate 
        localparam integer d727 = 27;
        for (n727 = 0; n727 < 16; n727 = n727 + 1) 
        begin: outbit727
            assign data_11[n727 + d727*16 + c25*28*16] = data_11_array[c25][d727][n727];
        end
    endgenerate
    localparam integer c26 = 26;
    generate 
        localparam integer d728 = 0;
        for (n728 = 0; n728 < 16; n728 = n728 + 1) 
        begin: outbit728
            assign data_11[n728 + d728*16 + c26*28*16] = data_11_array[c26][d728][n728];
        end
    endgenerate
    generate 
        localparam integer d729 = 1;
        for (n729 = 0; n729 < 16; n729 = n729 + 1) 
        begin: outbit729
            assign data_11[n729 + d729*16 + c26*28*16] = data_11_array[c26][d729][n729];
        end
    endgenerate
    generate 
        localparam integer d730 = 2;
        for (n730 = 0; n730 < 16; n730 = n730 + 1) 
        begin: outbit730
            assign data_11[n730 + d730*16 + c26*28*16] = data_11_array[c26][d730][n730];
        end
    endgenerate
    generate 
        localparam integer d731 = 3;
        for (n731 = 0; n731 < 16; n731 = n731 + 1) 
        begin: outbit731
            assign data_11[n731 + d731*16 + c26*28*16] = data_11_array[c26][d731][n731];
        end
    endgenerate
    generate 
        localparam integer d732 = 4;
        for (n732 = 0; n732 < 16; n732 = n732 + 1) 
        begin: outbit732
            assign data_11[n732 + d732*16 + c26*28*16] = data_11_array[c26][d732][n732];
        end
    endgenerate
    generate 
        localparam integer d733 = 5;
        for (n733 = 0; n733 < 16; n733 = n733 + 1) 
        begin: outbit733
            assign data_11[n733 + d733*16 + c26*28*16] = data_11_array[c26][d733][n733];
        end
    endgenerate
    generate 
        localparam integer d734 = 6;
        for (n734 = 0; n734 < 16; n734 = n734 + 1) 
        begin: outbit734
            assign data_11[n734 + d734*16 + c26*28*16] = data_11_array[c26][d734][n734];
        end
    endgenerate
    generate 
        localparam integer d735 = 7;
        for (n735 = 0; n735 < 16; n735 = n735 + 1) 
        begin: outbit735
            assign data_11[n735 + d735*16 + c26*28*16] = data_11_array[c26][d735][n735];
        end
    endgenerate
    generate 
        localparam integer d736 = 8;
        for (n736 = 0; n736 < 16; n736 = n736 + 1) 
        begin: outbit736
            assign data_11[n736 + d736*16 + c26*28*16] = data_11_array[c26][d736][n736];
        end
    endgenerate
    generate 
        localparam integer d737 = 9;
        for (n737 = 0; n737 < 16; n737 = n737 + 1) 
        begin: outbit737
            assign data_11[n737 + d737*16 + c26*28*16] = data_11_array[c26][d737][n737];
        end
    endgenerate
    generate 
        localparam integer d738 = 10;
        for (n738 = 0; n738 < 16; n738 = n738 + 1) 
        begin: outbit738
            assign data_11[n738 + d738*16 + c26*28*16] = data_11_array[c26][d738][n738];
        end
    endgenerate
    generate 
        localparam integer d739 = 11;
        for (n739 = 0; n739 < 16; n739 = n739 + 1) 
        begin: outbit739
            assign data_11[n739 + d739*16 + c26*28*16] = data_11_array[c26][d739][n739];
        end
    endgenerate
    generate 
        localparam integer d740 = 12;
        for (n740 = 0; n740 < 16; n740 = n740 + 1) 
        begin: outbit740
            assign data_11[n740 + d740*16 + c26*28*16] = data_11_array[c26][d740][n740];
        end
    endgenerate
    generate 
        localparam integer d741 = 13;
        for (n741 = 0; n741 < 16; n741 = n741 + 1) 
        begin: outbit741
            assign data_11[n741 + d741*16 + c26*28*16] = data_11_array[c26][d741][n741];
        end
    endgenerate
    generate 
        localparam integer d742 = 14;
        for (n742 = 0; n742 < 16; n742 = n742 + 1) 
        begin: outbit742
            assign data_11[n742 + d742*16 + c26*28*16] = data_11_array[c26][d742][n742];
        end
    endgenerate
    generate 
        localparam integer d743 = 15;
        for (n743 = 0; n743 < 16; n743 = n743 + 1) 
        begin: outbit743
            assign data_11[n743 + d743*16 + c26*28*16] = data_11_array[c26][d743][n743];
        end
    endgenerate
    generate 
        localparam integer d744 = 16;
        for (n744 = 0; n744 < 16; n744 = n744 + 1) 
        begin: outbit744
            assign data_11[n744 + d744*16 + c26*28*16] = data_11_array[c26][d744][n744];
        end
    endgenerate
    generate 
        localparam integer d745 = 17;
        for (n745 = 0; n745 < 16; n745 = n745 + 1) 
        begin: outbit745
            assign data_11[n745 + d745*16 + c26*28*16] = data_11_array[c26][d745][n745];
        end
    endgenerate
    generate 
        localparam integer d746 = 18;
        for (n746 = 0; n746 < 16; n746 = n746 + 1) 
        begin: outbit746
            assign data_11[n746 + d746*16 + c26*28*16] = data_11_array[c26][d746][n746];
        end
    endgenerate
    generate 
        localparam integer d747 = 19;
        for (n747 = 0; n747 < 16; n747 = n747 + 1) 
        begin: outbit747
            assign data_11[n747 + d747*16 + c26*28*16] = data_11_array[c26][d747][n747];
        end
    endgenerate
    generate 
        localparam integer d748 = 20;
        for (n748 = 0; n748 < 16; n748 = n748 + 1) 
        begin: outbit748
            assign data_11[n748 + d748*16 + c26*28*16] = data_11_array[c26][d748][n748];
        end
    endgenerate
    generate 
        localparam integer d749 = 21;
        for (n749 = 0; n749 < 16; n749 = n749 + 1) 
        begin: outbit749
            assign data_11[n749 + d749*16 + c26*28*16] = data_11_array[c26][d749][n749];
        end
    endgenerate
    generate 
        localparam integer d750 = 22;
        for (n750 = 0; n750 < 16; n750 = n750 + 1) 
        begin: outbit750
            assign data_11[n750 + d750*16 + c26*28*16] = data_11_array[c26][d750][n750];
        end
    endgenerate
    generate 
        localparam integer d751 = 23;
        for (n751 = 0; n751 < 16; n751 = n751 + 1) 
        begin: outbit751
            assign data_11[n751 + d751*16 + c26*28*16] = data_11_array[c26][d751][n751];
        end
    endgenerate
    generate 
        localparam integer d752 = 24;
        for (n752 = 0; n752 < 16; n752 = n752 + 1) 
        begin: outbit752
            assign data_11[n752 + d752*16 + c26*28*16] = data_11_array[c26][d752][n752];
        end
    endgenerate
    generate 
        localparam integer d753 = 25;
        for (n753 = 0; n753 < 16; n753 = n753 + 1) 
        begin: outbit753
            assign data_11[n753 + d753*16 + c26*28*16] = data_11_array[c26][d753][n753];
        end
    endgenerate
    generate 
        localparam integer d754 = 26;
        for (n754 = 0; n754 < 16; n754 = n754 + 1) 
        begin: outbit754
            assign data_11[n754 + d754*16 + c26*28*16] = data_11_array[c26][d754][n754];
        end
    endgenerate
    generate 
        localparam integer d755 = 27;
        for (n755 = 0; n755 < 16; n755 = n755 + 1) 
        begin: outbit755
            assign data_11[n755 + d755*16 + c26*28*16] = data_11_array[c26][d755][n755];
        end
    endgenerate
    localparam integer c27 = 27;
    generate 
        localparam integer d756 = 0;
        for (n756 = 0; n756 < 16; n756 = n756 + 1) 
        begin: outbit756
            assign data_11[n756 + d756*16 + c27*28*16] = data_11_array[c27][d756][n756];
        end
    endgenerate
    generate 
        localparam integer d757 = 1;
        for (n757 = 0; n757 < 16; n757 = n757 + 1) 
        begin: outbit757
            assign data_11[n757 + d757*16 + c27*28*16] = data_11_array[c27][d757][n757];
        end
    endgenerate
    generate 
        localparam integer d758 = 2;
        for (n758 = 0; n758 < 16; n758 = n758 + 1) 
        begin: outbit758
            assign data_11[n758 + d758*16 + c27*28*16] = data_11_array[c27][d758][n758];
        end
    endgenerate
    generate 
        localparam integer d759 = 3;
        for (n759 = 0; n759 < 16; n759 = n759 + 1) 
        begin: outbit759
            assign data_11[n759 + d759*16 + c27*28*16] = data_11_array[c27][d759][n759];
        end
    endgenerate
    generate 
        localparam integer d760 = 4;
        for (n760 = 0; n760 < 16; n760 = n760 + 1) 
        begin: outbit760
            assign data_11[n760 + d760*16 + c27*28*16] = data_11_array[c27][d760][n760];
        end
    endgenerate
    generate 
        localparam integer d761 = 5;
        for (n761 = 0; n761 < 16; n761 = n761 + 1) 
        begin: outbit761
            assign data_11[n761 + d761*16 + c27*28*16] = data_11_array[c27][d761][n761];
        end
    endgenerate
    generate 
        localparam integer d762 = 6;
        for (n762 = 0; n762 < 16; n762 = n762 + 1) 
        begin: outbit762
            assign data_11[n762 + d762*16 + c27*28*16] = data_11_array[c27][d762][n762];
        end
    endgenerate
    generate 
        localparam integer d763 = 7;
        for (n763 = 0; n763 < 16; n763 = n763 + 1) 
        begin: outbit763
            assign data_11[n763 + d763*16 + c27*28*16] = data_11_array[c27][d763][n763];
        end
    endgenerate
    generate 
        localparam integer d764 = 8;
        for (n764 = 0; n764 < 16; n764 = n764 + 1) 
        begin: outbit764
            assign data_11[n764 + d764*16 + c27*28*16] = data_11_array[c27][d764][n764];
        end
    endgenerate
    generate 
        localparam integer d765 = 9;
        for (n765 = 0; n765 < 16; n765 = n765 + 1) 
        begin: outbit765
            assign data_11[n765 + d765*16 + c27*28*16] = data_11_array[c27][d765][n765];
        end
    endgenerate
    generate 
        localparam integer d766 = 10;
        for (n766 = 0; n766 < 16; n766 = n766 + 1) 
        begin: outbit766
            assign data_11[n766 + d766*16 + c27*28*16] = data_11_array[c27][d766][n766];
        end
    endgenerate
    generate 
        localparam integer d767 = 11;
        for (n767 = 0; n767 < 16; n767 = n767 + 1) 
        begin: outbit767
            assign data_11[n767 + d767*16 + c27*28*16] = data_11_array[c27][d767][n767];
        end
    endgenerate
    generate 
        localparam integer d768 = 12;
        for (n768 = 0; n768 < 16; n768 = n768 + 1) 
        begin: outbit768
            assign data_11[n768 + d768*16 + c27*28*16] = data_11_array[c27][d768][n768];
        end
    endgenerate
    generate 
        localparam integer d769 = 13;
        for (n769 = 0; n769 < 16; n769 = n769 + 1) 
        begin: outbit769
            assign data_11[n769 + d769*16 + c27*28*16] = data_11_array[c27][d769][n769];
        end
    endgenerate
    generate 
        localparam integer d770 = 14;
        for (n770 = 0; n770 < 16; n770 = n770 + 1) 
        begin: outbit770
            assign data_11[n770 + d770*16 + c27*28*16] = data_11_array[c27][d770][n770];
        end
    endgenerate
    generate 
        localparam integer d771 = 15;
        for (n771 = 0; n771 < 16; n771 = n771 + 1) 
        begin: outbit771
            assign data_11[n771 + d771*16 + c27*28*16] = data_11_array[c27][d771][n771];
        end
    endgenerate
    generate 
        localparam integer d772 = 16;
        for (n772 = 0; n772 < 16; n772 = n772 + 1) 
        begin: outbit772
            assign data_11[n772 + d772*16 + c27*28*16] = data_11_array[c27][d772][n772];
        end
    endgenerate
    generate 
        localparam integer d773 = 17;
        for (n773 = 0; n773 < 16; n773 = n773 + 1) 
        begin: outbit773
            assign data_11[n773 + d773*16 + c27*28*16] = data_11_array[c27][d773][n773];
        end
    endgenerate
    generate 
        localparam integer d774 = 18;
        for (n774 = 0; n774 < 16; n774 = n774 + 1) 
        begin: outbit774
            assign data_11[n774 + d774*16 + c27*28*16] = data_11_array[c27][d774][n774];
        end
    endgenerate
    generate 
        localparam integer d775 = 19;
        for (n775 = 0; n775 < 16; n775 = n775 + 1) 
        begin: outbit775
            assign data_11[n775 + d775*16 + c27*28*16] = data_11_array[c27][d775][n775];
        end
    endgenerate
    generate 
        localparam integer d776 = 20;
        for (n776 = 0; n776 < 16; n776 = n776 + 1) 
        begin: outbit776
            assign data_11[n776 + d776*16 + c27*28*16] = data_11_array[c27][d776][n776];
        end
    endgenerate
    generate 
        localparam integer d777 = 21;
        for (n777 = 0; n777 < 16; n777 = n777 + 1) 
        begin: outbit777
            assign data_11[n777 + d777*16 + c27*28*16] = data_11_array[c27][d777][n777];
        end
    endgenerate
    generate 
        localparam integer d778 = 22;
        for (n778 = 0; n778 < 16; n778 = n778 + 1) 
        begin: outbit778
            assign data_11[n778 + d778*16 + c27*28*16] = data_11_array[c27][d778][n778];
        end
    endgenerate
    generate 
        localparam integer d779 = 23;
        for (n779 = 0; n779 < 16; n779 = n779 + 1) 
        begin: outbit779
            assign data_11[n779 + d779*16 + c27*28*16] = data_11_array[c27][d779][n779];
        end
    endgenerate
    generate 
        localparam integer d780 = 24;
        for (n780 = 0; n780 < 16; n780 = n780 + 1) 
        begin: outbit780
            assign data_11[n780 + d780*16 + c27*28*16] = data_11_array[c27][d780][n780];
        end
    endgenerate
    generate 
        localparam integer d781 = 25;
        for (n781 = 0; n781 < 16; n781 = n781 + 1) 
        begin: outbit781
            assign data_11[n781 + d781*16 + c27*28*16] = data_11_array[c27][d781][n781];
        end
    endgenerate
    generate 
        localparam integer d782 = 26;
        for (n782 = 0; n782 < 16; n782 = n782 + 1) 
        begin: outbit782
            assign data_11[n782 + d782*16 + c27*28*16] = data_11_array[c27][d782][n782];
        end
    endgenerate
    generate 
        localparam integer d783 = 27;
        for (n783 = 0; n783 < 16; n783 = n783 + 1) 
        begin: outbit783
            assign data_11[n783 + d783*16 + c27*28*16] = data_11_array[c27][d783][n783];
        end
    endgenerate

endmodule
